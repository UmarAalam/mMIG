// Benchmark "metricComp" written by ABC on Wed Apr 29 17:58:01 2015

module metricComp ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192;
  wire n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
    n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
    n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
    n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
    n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
    n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
    n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
    n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
    n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
    n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
    n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
    n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
    n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
    n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5746, n5747,
    n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
    n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
    n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
    n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
    n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
    n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
    n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
    n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
    n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
    n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
    n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
    n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
    n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
    n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
    n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
    n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
    n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
    n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
    n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
    n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
    n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
    n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
    n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
    n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
    n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
    n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
    n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
    n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
    n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
    n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
    n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6718,
    n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
    n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
    n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
    n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
    n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
    n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
    n8962, n8963, n8964, n8965, n8966, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
    n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
    n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
    n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
    n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
    n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
    n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
    n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
    n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
    n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
    n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
    n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
    n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
    n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
    n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
    n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
    n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
    n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
    n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
    n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
    n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
    n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
    n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
    n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
    n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
    n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
    n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
    n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
    n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
    n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
    n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
    n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
    n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
    n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
    n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
    n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
    n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
    n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
    n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
    n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
    n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
    n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
    n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
    n11472, n11473, n11474, n11475, n11476, n11478, n11479, n11480, n11481,
    n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
    n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
    n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
    n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
    n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
    n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
    n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
    n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
    n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
    n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
    n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
    n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
    n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
    n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
    n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
    n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
    n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
    n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
    n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
    n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
    n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
    n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
    n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
    n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
    n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
    n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
    n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
    n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
    n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
    n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
    n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
    n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
    n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
    n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
    n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
    n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
    n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
    n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
    n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
    n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
    n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
    n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
    n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
    n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
    n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
    n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
    n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
    n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
    n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
    n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
    n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
    n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
    n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
    n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
    n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
    n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
    n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
    n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
    n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
    n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
    n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
    n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
    n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
    n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
    n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
    n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
    n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
    n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
    n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
    n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
    n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
    n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
    n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
    n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
    n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
    n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
    n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
    n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
    n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
    n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
    n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
    n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
    n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
    n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
    n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
    n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
    n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
    n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
    n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
    n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
    n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
    n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
    n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
    n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
    n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
    n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
    n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
    n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
    n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
    n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
    n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
    n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
    n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
    n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
    n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
    n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
    n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
    n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
    n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
    n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
    n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
    n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
    n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
    n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
    n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
    n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
    n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
    n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
    n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
    n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
    n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
    n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
    n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
    n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
    n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
    n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
    n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
    n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
    n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
    n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
    n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
    n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
    n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
    n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
    n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
    n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
    n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
    n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
    n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
    n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
    n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
    n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
    n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
    n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
    n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
    n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
    n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
    n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
    n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
    n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
    n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
    n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
    n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
    n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
    n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
    n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
    n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
    n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
    n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
    n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
    n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
    n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
    n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
    n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
    n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
    n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
    n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
    n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
    n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
    n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
    n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16208, n16209,
    n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
    n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
    n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
    n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
    n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
    n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
    n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
    n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
    n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
    n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
    n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
    n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
    n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
    n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
    n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
    n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
    n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
    n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
    n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
    n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
    n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
    n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
    n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
    n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
    n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
    n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
    n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
    n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
    n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
    n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
    n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
    n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
    n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
    n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
    n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
    n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
    n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
    n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
    n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
    n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
    n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
    n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
    n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
    n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
    n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
    n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
    n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
    n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
    n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
    n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
    n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
    n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
    n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
    n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
    n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
    n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
    n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
    n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
    n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
    n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
    n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
    n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
    n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
    n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
    n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
    n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
    n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
    n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
    n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
    n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
    n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
    n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
    n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
    n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
    n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
    n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
    n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
    n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
    n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
    n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
    n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
    n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
    n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
    n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
    n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
    n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
    n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
    n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
    n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
    n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
    n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
    n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
    n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
    n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
    n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
    n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
    n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
    n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
    n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
    n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
    n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
    n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
    n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
    n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
    n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
    n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
    n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
    n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
    n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
    n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
    n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
    n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
    n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
    n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
    n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
    n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
    n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
    n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
    n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
    n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
    n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
    n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
    n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
    n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
    n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
    n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
    n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
    n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
    n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
    n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
    n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
    n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
    n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
    n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
    n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
    n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
    n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
    n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
    n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
    n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
    n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
    n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
    n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
    n18174, n18175, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199, n18201, n18202, n18203,
    n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
    n18223, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
    n18233, n18234, n18235, n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18249, n18250, n18251, n18252,
    n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
    n18271, n18272, n18273, n18274, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
    n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
    n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18411,
    n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
    n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
    n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18503, n18504,
    n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
    n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
    n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
    n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
    n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
    n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18731, n18732, n18733, n18734, n18735,
    n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
    n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
    n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
    n18763, n18764, n18765, n18766, n18767, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
    n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18887, n18888, n18889, n18890, n18891,
    n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
    n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
    n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
    n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
    n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
    n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
    n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
    n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19064, n19065,
    n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
    n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
    n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
    n19120, n19121, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
    n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
    n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
    n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
    n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
    n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
    n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
    n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
    n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
    n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
    n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
    n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
    n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
    n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19473, n19474, n19475, n19476,
    n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
    n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
    n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
    n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
    n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
    n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
    n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
    n19540, n19541, n19542, n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
    n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
    n19613, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
    n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
    n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
    n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19686,
    n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
    n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
    n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
    n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
    n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
    n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
    n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
    n19750, n19751, n19752, n19753, n19754, n19755, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
    n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
    n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
    n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
    n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19938, n19939, n19940, n19941,
    n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
    n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
    n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
    n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
    n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
    n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
    n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
    n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
    n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
    n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
    n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
    n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
    n20141, n20142, n20143, n20144, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
    n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
    n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
    n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
    n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
    n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
    n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
    n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
    n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
    n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
    n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
    n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
    n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
    n20350, n20351, n20352, n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
    n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
    n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20458, n20459,
    n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
    n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
    n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
    n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
    n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
    n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
    n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
    n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
    n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
    n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
    n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
    n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
    n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
    n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
    n20659, n20660, n20661, n20662, n20663, n20664, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20813,
    n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
    n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
    n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
    n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
    n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20939, n20940,
    n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
    n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
    n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
    n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
    n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
    n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
    n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
    n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
    n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
    n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
    n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
    n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
    n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
    n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21189, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
    n21312, n21313, n21314, n21315, n21317, n21318, n21319, n21320, n21321,
    n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
    n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
    n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
    n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
    n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
    n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
    n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
    n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
    n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
    n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
    n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
    n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
    n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
    n21439, n21440, n21441, n21443, n21444, n21445, n21446, n21447, n21448,
    n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
    n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
    n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
    n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
    n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
    n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
    n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
    n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
    n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
    n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
    n21566, n21567, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
    n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
    n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
    n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
    n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
    n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
    n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
    n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
    n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
    n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
    n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
    n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
    n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
    n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
    n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
    n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
    n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
    n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
    n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
    n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
    n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
    n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
    n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
    n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
    n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
    n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
    n21865, n21866, n21867, n21868, n21869, n21870, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
    n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
    n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
    n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
    n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
    n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
    n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
    n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
    n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
    n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
    n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
    n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
    n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22203, n22204, n22206, n22207, n22208, n22209,
    n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
    n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
    n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
    n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
    n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
    n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
    n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
    n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
    n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
    n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
    n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
    n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
    n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
    n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
    n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
    n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22707,
    n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
    n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
    n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
    n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
    n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
    n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
    n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
    n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
    n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
    n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
    n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
    n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
    n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
    n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
    n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
    n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
    n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
    n22870, n22871, n22872, n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
    n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
    n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
    n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
    n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
    n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
    n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
    n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
    n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
    n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
    n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
    n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
    n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
    n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
    n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
    n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
    n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
    n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
    n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
    n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
    n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
    n23250, n23251, n23252, n23253, n23255, n23256, n23257, n23258, n23259,
    n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
    n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
    n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
    n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
    n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
    n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
    n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
    n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
    n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
    n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
    n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
    n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
    n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
    n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
    n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
    n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
    n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
    n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
    n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
    n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
    n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
    n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
    n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
    n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
    n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
    n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
    n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
    n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
    n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
    n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
    n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
    n23639, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
    n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
    n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
    n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
    n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
    n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
    n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
    n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
    n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
    n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
    n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23834, n23835, n23836, n23837, n23838,
    n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
    n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
    n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
    n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
    n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
    n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
    n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910,
    n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
    n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
    n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
    n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
    n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
    n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
    n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
    n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982,
    n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
    n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
    n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
    n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
    n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
    n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
    n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
    n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
    n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
    n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24413, n24414, n24415, n24416, n24417,
    n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
    n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
    n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
    n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462,
    n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
    n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
    n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
    n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
    n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
    n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516,
    n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
    n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
    n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
    n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
    n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
    n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
    n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
    n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588,
    n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
    n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847, n24849, n24850, n24851,
    n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
    n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869,
    n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
    n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
    n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
    n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
    n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
    n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
    n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
    n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941,
    n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950,
    n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
    n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
    n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
    n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
    n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
    n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
    n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
    n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
    n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
    n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
    n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
    n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
    n25077, n25078, n25079, n25080, n25082, n25083, n25084, n25085, n25086,
    n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
    n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
    n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
    n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
    n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
    n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140,
    n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
    n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
    n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
    n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
    n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
    n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
    n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
    n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212,
    n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
    n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230,
    n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
    n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
    n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
    n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
    n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
    n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284,
    n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
    n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
    n25312, n25313, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
    n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
    n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
    n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
    n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
    n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
    n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
    n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
    n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
    n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
    n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
    n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
    n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
    n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
    n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
    n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
    n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
    n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
    n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
    n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
    n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
    n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
    n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
    n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
    n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
    n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
    n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
    n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
    n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25781, n25782,
    n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
    n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
    n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
    n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
    n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
    n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
    n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
    n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
    n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
    n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
    n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
    n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
    n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
    n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
    n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
    n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
    n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
    n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
    n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
    n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
    n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
    n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
    n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
    n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
    n26008, n26009, n26010, n26011, n26012, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
    n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
    n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
    n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
    n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
    n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
    n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
    n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
    n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
    n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
    n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
    n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
    n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
    n26243, n26244, n26245, n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
    n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
    n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
    n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
    n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
    n26478, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
    n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
    n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
    n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
    n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
    n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
    n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541,
    n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550,
    n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
    n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
    n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
    n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
    n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
    n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
    n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
    n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
    n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
    n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
    n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
    n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
    n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
    n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
    n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
    n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694,
    n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
    n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
    n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
    n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
    n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
    n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
    n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
    n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766,
    n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
    n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
    n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
    n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
    n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
    n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
    n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
    n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27043, n27044, n27045, n27046, n27047,
    n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
    n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
    n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
    n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
    n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
    n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
    n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
    n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
    n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
    n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
    n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
    n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
    n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
    n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
    n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
    n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
    n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
    n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
    n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
    n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
    n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
    n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
    n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
    n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
    n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
    n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
    n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
    n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
    n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27309,
    n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
    n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
    n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
    n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
    n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
    n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
    n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
    n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381,
    n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390,
    n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
    n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
    n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
    n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
    n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
    n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
    n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453,
    n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
    n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
    n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
    n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
    n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
    n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
    n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
    n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
    n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534,
    n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543,
    n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
    n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
    n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
    n27571, n27572, n27573, n27575, n27576, n27577, n27578, n27579, n27580,
    n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
    n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
    n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
    n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
    n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
    n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
    n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
    n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
    n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832,
    n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
    n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
    n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
    n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
    n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
    n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
    n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
    n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
    n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
    n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
    n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
    n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
    n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
    n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
    n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
    n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
    n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
    n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
    n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
    n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
    n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
    n28104, n28105, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
    n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
    n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
    n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
    n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
    n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
    n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
    n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176,
    n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
    n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
    n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
    n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
    n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
    n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
    n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
    n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
    n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
    n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
    n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
    n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
    n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
    n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
    n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
    n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
    n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
    n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
    n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
    n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
    n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
    n28366, n28367, n28368, n28369, n28370, n28371, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
    n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
    n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
    n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
    n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
    n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
    n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
    n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
    n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
    n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
    n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
    n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
    n28637, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
    n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
    n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
    n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
    n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
    n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
    n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
    n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
    n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
    n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
    n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
    n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
    n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
    n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
    n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28972, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
    n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
    n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
    n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
    n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061,
    n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
    n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
    n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
    n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
    n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
    n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
    n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
    n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
    n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
    n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
    n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
    n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
    n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
    n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
    n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196,
    n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
    n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
    n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
    n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
    n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
    n29269, n29270, n29271, n29272, n29273, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29576,
    n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
    n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
    n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
    n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621,
    n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
    n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639,
    n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648,
    n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
    n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
    n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
    n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684,
    n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693,
    n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
    n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711,
    n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
    n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
    n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
    n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
    n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756,
    n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765,
    n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
    n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
    n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
    n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
    n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
    n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
    n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828,
    n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837,
    n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
    n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855,
    n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
    n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
    n29874, n29875, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
    n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892,
    n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901,
    n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
    n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
    n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
    n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
    n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
    n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
    n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964,
    n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973,
    n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
    n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
    n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
    n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
    n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
    n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
    n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036,
    n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045,
    n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
    n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
    n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
    n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
    n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
    n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
    n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
    n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117,
    n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
    n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135,
    n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
    n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
    n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
    n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
    n30172, n30173, n30174, n30175, n30176, n30178, n30179, n30180, n30181,
    n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
    n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
    n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
    n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
    n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
    n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
    n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244,
    n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253,
    n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
    n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
    n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
    n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
    n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
    n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
    n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
    n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388,
    n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397,
    n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
    n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
    n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
    n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
    n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
    n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
    n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
    n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469,
    n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30479,
    n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
    n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
    n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
    n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
    n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
    n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533,
    n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
    n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
    n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
    n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
    n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
    n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605,
    n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
    n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
    n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
    n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
    n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
    n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
    n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677,
    n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
    n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
    n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
    n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
    n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
    n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
    n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740,
    n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749,
    n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
    n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
    n30777, n30778, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
    n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
    n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804,
    n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813,
    n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
    n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
    n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
    n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
    n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
    n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
    n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876,
    n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885,
    n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
    n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
    n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
    n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
    n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
    n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
    n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948,
    n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957,
    n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
    n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
    n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
    n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
    n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
    n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
    n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020,
    n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029,
    n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
    n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
    n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
    n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
    n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074,
    n31075, n31076, n31077, n31078, n31079, n31081, n31082, n31083, n31084,
    n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
    n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
    n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
    n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
    n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
    n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
    n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
    n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
    n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
    n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
    n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
    n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
    n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
    n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
    n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
    n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
    n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
    n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381,
    n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
    n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
    n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
    n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
    n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
    n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
    n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453,
    n31454, n31455, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
    n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
    n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
    n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517,
    n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
    n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
    n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
    n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
    n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589,
    n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
    n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
    n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
    n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661,
    n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
    n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
    n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
    n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
    n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
    n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
    n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733,
    n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
    n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
    n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
    n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797,
    n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
    n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
    n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824,
    n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
    n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
    n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
    n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
    n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869,
    n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
    n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
    n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896,
    n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
    n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
    n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
    n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
    n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941,
    n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
    n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
    n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
    n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
    n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
    n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
    n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
    n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013,
    n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
    n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031,
    n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
    n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
    n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
    n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
    n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
    n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085,
    n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
    n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103,
    n32104, n32105, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
    n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
    n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149,
    n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
    n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
    n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
    n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
    n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
    n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
    n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
    n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
    n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
    n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
    n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
    n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
    n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
    n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
    n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
    n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
    n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
    n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
    n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
    n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
    n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
    n32429, n32430, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
    n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
    n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501,
    n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
    n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519,
    n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
    n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
    n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
    n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
    n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573,
    n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
    n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591,
    n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
    n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
    n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
    n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
    n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
    n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
    n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
    n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
    n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
    n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
    n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
    n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
    n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717,
    n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
    n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
    n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
    n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
    n32754, n32755, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
    n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772,
    n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781,
    n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
    n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799,
    n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808,
    n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
    n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
    n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
    n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844,
    n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853,
    n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
    n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871,
    n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880,
    n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
    n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
    n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
    n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916,
    n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925,
    n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
    n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
    n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
    n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
    n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
    n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
    n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997,
    n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
    n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
    n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024,
    n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
    n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
    n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
    n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069,
    n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
    n33079, n33080, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
    n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
    n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
    n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133,
    n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
    n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
    n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
    n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
    n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
    n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
    n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
    n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
    n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
    n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
    n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
    n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
    n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
    n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
    n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
    n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
    n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
    n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431,
    n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
    n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
    n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
    n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
    n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
    n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485,
    n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
    n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503,
    n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
    n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
    n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
    n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
    n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
    n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557,
    n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
    n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575,
    n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
    n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
    n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
    n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
    n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
    n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
    n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
    n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647,
    n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
    n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
    n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
    n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
    n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
    n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701,
    n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
    n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719,
    n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
    n33729, n33730, n33732, n33733, n33734, n33735, n33736, n33737, n33738,
    n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
    n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756,
    n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765,
    n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
    n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783,
    n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792,
    n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
    n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810,
    n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
    n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828,
    n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837,
    n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
    n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855,
    n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864,
    n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
    n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
    n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
    n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909,
    n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
    n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927,
    n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936,
    n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
    n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954,
    n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
    n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972,
    n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981,
    n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
    n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999,
    n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
    n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
    n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026,
    n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
    n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044,
    n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053,
    n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
    n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
    n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080,
    n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
    n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
    n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
    n34108, n34109, n34111, n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
    n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
    n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
    n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
    n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189,
    n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
    n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
    n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
    n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
    n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
    n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
    n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
    n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261,
    n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
    n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
    n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
    n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
    n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
    n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
    n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
    n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333,
    n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
    n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
    n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
    n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
    n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
    n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
    n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
    n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405,
    n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
    n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
    n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
    n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
    n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
    n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
    n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34483, n34484, n34485, n34486, n34487,
    n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
    n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
    n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
    n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
    n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
    n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541,
    n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
    n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
    n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
    n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
    n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
    n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
    n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
    n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613,
    n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
    n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
    n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
    n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
    n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
    n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
    n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685,
    n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
    n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
    n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
    n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
    n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
    n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
    n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757,
    n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
    n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
    n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
    n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
    n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
    n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
    n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
    n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829,
    n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
    n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
    n34848, n34849, n34850, n34851, n34852, n34853, n34855, n34856, n34857,
    n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
    n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
    n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884,
    n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893,
    n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
    n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911,
    n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920,
    n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
    n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
    n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
    n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956,
    n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965,
    n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
    n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983,
    n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992,
    n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
    n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010,
    n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
    n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028,
    n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037,
    n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
    n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055,
    n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064,
    n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
    n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082,
    n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
    n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100,
    n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109,
    n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
    n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
    n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
    n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
    n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154,
    n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
    n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172,
    n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181,
    n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
    n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199,
    n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208,
    n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
    n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
    n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
    n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
    n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
    n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
    n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
    n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
    n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
    n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
    n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
    n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
    n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
    n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
    n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
    n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
    n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
    n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
    n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
    n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
    n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
    n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
    n35597, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
    n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
    n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624,
    n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
    n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642,
    n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
    n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660,
    n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669,
    n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
    n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687,
    n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696,
    n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
    n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714,
    n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
    n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732,
    n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741,
    n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
    n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
    n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768,
    n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
    n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
    n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
    n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813,
    n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
    n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831,
    n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840,
    n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
    n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858,
    n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
    n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885,
    n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
    n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
    n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
    n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
    n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
    n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948,
    n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957,
    n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
    n35967, n35968, n35969, n35971, n35972, n35973, n35974, n35975, n35976,
    n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
    n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
    n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
    n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012,
    n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021,
    n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
    n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
    n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048,
    n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
    n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
    n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
    n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084,
    n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093,
    n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
    n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111,
    n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
    n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
    n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138,
    n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
    n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156,
    n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165,
    n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
    n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183,
    n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
    n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
    n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210,
    n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
    n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228,
    n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237,
    n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
    n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255,
    n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264,
    n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
    n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282,
    n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
    n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300,
    n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309,
    n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
    n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327,
    n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336,
    n36337, n36338, n36339, n36340, n36341, n36343, n36344, n36345, n36346,
    n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
    n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364,
    n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
    n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400,
    n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
    n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436,
    n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445,
    n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
    n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
    n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
    n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508,
    n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
    n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
    n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
    n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
    n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580,
    n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589,
    n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
    n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
    n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616,
    n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
    n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
    n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
    n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652,
    n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661,
    n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
    n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679,
    n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688,
    n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
    n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
    n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36715, n36716,
    n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725,
    n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
    n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
    n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752,
    n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
    n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
    n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
    n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788,
    n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797,
    n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
    n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815,
    n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824,
    n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
    n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
    n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860,
    n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869,
    n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
    n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887,
    n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
    n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
    n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
    n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
    n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932,
    n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941,
    n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
    n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
    n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
    n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
    n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
    n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
    n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004,
    n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013,
    n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031,
    n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
    n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
    n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
    n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
    n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076,
    n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085,
    n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
    n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103,
    n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
    n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
    n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140,
    n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149,
    n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
    n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167,
    n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176,
    n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
    n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
    n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
    n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212,
    n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221,
    n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
    n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239,
    n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248,
    n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
    n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
    n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
    n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284,
    n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293,
    n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
    n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311,
    n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320,
    n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
    n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
    n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
    n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356,
    n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365,
    n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
    n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383,
    n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
    n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
    n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
    n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
    n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428,
    n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437,
    n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
    n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455,
    n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
    n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
    n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
    n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
    n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
    n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
    n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
    n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
    n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
    n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573,
    n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
    n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
    n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
    n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
    n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
    n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
    n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
    n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
    n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
    n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
    n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708,
    n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717,
    n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
    n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735,
    n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
    n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
    n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
    n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
    n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780,
    n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789,
    n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
    n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807,
    n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
    n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
    n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
    n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
    n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852,
    n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861,
    n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
    n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879,
    n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
    n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
    n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
    n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
    n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924,
    n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933,
    n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
    n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
    n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
    n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
    n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
    n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997,
    n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
    n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
    n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
    n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
    n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
    n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
    n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
    n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
    n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
    n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
    n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
    n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
    n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
    n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
    n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204,
    n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
    n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
    n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276,
    n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285,
    n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
    n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
    n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
    n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
    n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349,
    n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
    n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367,
    n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376,
    n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
    n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
    n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403,
    n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412,
    n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421,
    n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
    n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439,
    n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
    n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
    n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
    n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
    n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484,
    n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493,
    n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
    n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511,
    n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
    n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
    n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
    n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
    n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556,
    n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565,
    n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
    n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583,
    n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
    n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
    n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
    n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
    n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628,
    n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637,
    n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
    n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655,
    n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
    n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
    n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
    n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691,
    n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700,
    n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709,
    n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
    n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727,
    n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
    n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
    n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
    n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764,
    n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
    n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
    n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
    n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
    n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
    n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836,
    n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845,
    n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
    n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
    n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
    n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
    n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
    n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
    n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
    n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917,
    n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
    n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
    n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
    n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989,
    n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
    n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
    n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
    n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
    n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052,
    n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
    n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
    n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
    n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124,
    n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
    n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
    n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
    n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
    n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
    n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188,
    n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197,
    n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
    n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215,
    n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
    n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
    n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
    n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
    n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260,
    n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269,
    n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
    n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
    n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
    n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
    n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
    n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
    n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332,
    n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341,
    n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
    n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359,
    n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
    n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
    n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
    n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395,
    n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404,
    n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413,
    n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
    n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431,
    n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
    n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
    n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
    n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467,
    n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476,
    n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484, n39485,
    n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494,
    n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503,
    n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
    n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
    n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
    n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
    n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548,
    n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557,
    n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567,
    n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
    n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
    n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
    n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
    n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612,
    n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621,
    n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630,
    n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639,
    n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
    n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
    n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
    n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675,
    n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684,
    n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693,
    n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702,
    n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711,
    n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
    n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
    n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
    n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747,
    n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756,
    n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764, n39765,
    n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
    n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783,
    n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
    n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
    n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
    n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
    n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828,
    n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837,
    n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
    n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855,
    n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
    n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
    n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
    n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891,
    n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900,
    n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908, n39909,
    n39910, n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
    n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927,
    n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
    n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
    n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
    n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963,
    n39966, n39968, n39970, n39971, n39973, n39975, n39977, n39978, n39979,
    n39981, n39982, n39984, n39985, n39986, n39988, n39989, n39990, n39991,
    n39993, n39994, n39995, n39996, n39998, n39999, n40000, n40001, n40002,
    n40004, n40005, n40006, n40007, n40008, n40009, n40011, n40012, n40013,
    n40014, n40015, n40017, n40018, n40019, n40020, n40021, n40022, n40024,
    n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40033, n40034,
    n40035, n40036, n40037, n40038, n40039, n40040, n40042, n40043, n40044,
    n40045, n40046, n40047, n40048, n40050, n40051, n40052, n40053, n40054,
    n40055, n40056, n40057, n40059, n40060, n40061, n40062, n40063, n40064,
    n40065, n40066, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
    n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084,
    n40085, n40086, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
    n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
    n40115, n40116, n40117, n40118, n40120, n40121, n40122, n40123, n40124,
    n40125, n40126, n40127, n40128, n40129, n40131, n40132, n40133, n40134,
    n40135, n40136, n40137, n40139, n40140, n40141, n40142, n40143, n40144,
    n40145, n40146, n40147, n40148, n40149, n40151, n40152, n40153, n40154,
    n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40163, n40164,
    n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173,
    n40174, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183,
    n40184, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
    n40194, n40195, n40196, n40197, n40198, n40199, n40201, n40202, n40203,
    n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212,
    n40213, n40214, n40215, n40217, n40218, n40219, n40220, n40221, n40222,
    n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
    n40242, n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251,
    n40252, n40253, n40254, n40255, n40256, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
    n40271, n40272, n40273, n40274, n40275, n40277, n40278, n40279, n40280,
    n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
    n40290, n40291, n40292, n40293, n40294, n40295, n40297, n40298, n40299,
    n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308,
    n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317,
    n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
    n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335,
    n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
    n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
    n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
    n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371,
    n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380,
    n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389,
    n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
    n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407,
    n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
    n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
    n40426, n40427, n40428, n40430, n40431, n40432, n40433, n40434, n40435,
    n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444,
    n40445, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
    n40464, n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
    n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
    n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
    n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500,
    n40501, n40502, n40503, n40504, n40505, n40506;
  assign n473 = ~pi042 & pi050;
  assign n474 = pi042 & ~pi050;
  assign n475 = ~pi043 & pi051;
  assign n476 = pi043 & ~pi051;
  assign n477 = ~pi044 & pi052;
  assign n478 = pi044 & ~pi052;
  assign n479 = pi046 & ~pi054;
  assign n480 = pi045 & ~pi053;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~pi045 & pi053;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n478 & ~n483;
  assign n485 = ~n477 & ~n484;
  assign n486 = ~n476 & ~n485;
  assign n487 = ~n475 & ~n486;
  assign n488 = ~n474 & ~n487;
  assign n489 = ~n473 & ~n488;
  assign n490 = ~pi041 & ~n489;
  assign n491 = pi041 & ~n473;
  assign n492 = ~n488 & n491;
  assign n493 = pi049 & ~n492;
  assign n494 = ~pi040 & pi048;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n490 & n495;
  assign n497 = pi040 & ~pi048;
  assign n498 = pi039 & ~pi047;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n496 & n499;
  assign n501 = ~pi039 & pi047;
  assign n502 = pi002 & ~n501;
  assign n503 = ~n500 & n502;
  assign n504 = ~pi039 & pi079;
  assign n505 = ~pi042 & pi082;
  assign n506 = pi042 & ~pi082;
  assign n507 = ~pi043 & pi083;
  assign n508 = pi043 & ~pi083;
  assign n509 = ~pi044 & pi084;
  assign n510 = pi044 & ~pi084;
  assign n511 = pi046 & ~pi086;
  assign n512 = pi045 & ~pi085;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~pi045 & pi085;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n510 & ~n515;
  assign n517 = ~n509 & ~n516;
  assign n518 = ~n508 & ~n517;
  assign n519 = ~n507 & ~n518;
  assign n520 = ~n506 & ~n519;
  assign n521 = ~n505 & ~n520;
  assign n522 = ~pi041 & ~n521;
  assign n523 = pi041 & ~n505;
  assign n524 = ~n520 & n523;
  assign n525 = pi081 & ~n524;
  assign n526 = ~pi040 & pi080;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~n522 & n527;
  assign n529 = pi040 & ~pi080;
  assign n530 = pi039 & ~pi079;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n528 & n531;
  assign n533 = ~n504 & ~n532;
  assign n534 = ~pi039 & pi095;
  assign n535 = ~pi042 & pi098;
  assign n536 = pi042 & ~pi098;
  assign n537 = ~pi043 & pi099;
  assign n538 = pi043 & ~pi099;
  assign n539 = ~pi044 & pi100;
  assign n540 = pi044 & ~pi100;
  assign n541 = pi046 & ~pi102;
  assign n542 = pi045 & ~pi101;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~pi045 & pi101;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n540 & ~n545;
  assign n547 = ~n539 & ~n546;
  assign n548 = ~n538 & ~n547;
  assign n549 = ~n537 & ~n548;
  assign n550 = ~n536 & ~n549;
  assign n551 = ~n535 & ~n550;
  assign n552 = ~pi041 & ~n551;
  assign n553 = pi041 & ~n535;
  assign n554 = ~n550 & n553;
  assign n555 = pi097 & ~n554;
  assign n556 = ~pi040 & pi096;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~n552 & n557;
  assign n559 = pi040 & ~pi096;
  assign n560 = pi039 & ~pi095;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n558 & n561;
  assign n563 = ~n534 & ~n562;
  assign n564 = ~n533 & ~n563;
  assign po144 = ~n500 & ~n501;
  assign n566 = ~pi039 & pi063;
  assign n567 = ~pi042 & pi066;
  assign n568 = pi042 & ~pi066;
  assign n569 = ~pi043 & pi067;
  assign n570 = pi043 & ~pi067;
  assign n571 = ~pi044 & pi068;
  assign n572 = pi044 & ~pi068;
  assign n573 = pi046 & ~pi070;
  assign n574 = pi045 & ~pi069;
  assign n575 = ~n573 & ~n574;
  assign n576 = ~pi045 & pi069;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~n572 & ~n577;
  assign n579 = ~n571 & ~n578;
  assign n580 = ~n570 & ~n579;
  assign n581 = ~n569 & ~n580;
  assign n582 = ~n568 & ~n581;
  assign n583 = ~n567 & ~n582;
  assign n584 = ~pi041 & ~n583;
  assign n585 = pi041 & ~n567;
  assign n586 = ~n582 & n585;
  assign n587 = pi065 & ~n586;
  assign n588 = ~pi040 & pi064;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n584 & n589;
  assign n591 = pi040 & ~pi064;
  assign n592 = pi039 & ~pi063;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n590 & n593;
  assign n595 = ~n566 & ~n594;
  assign n596 = ~po144 & ~n595;
  assign n597 = n564 & n596;
  assign n598 = ~pi039 & pi199;
  assign n599 = ~pi042 & pi202;
  assign n600 = pi042 & ~pi202;
  assign n601 = ~pi043 & pi203;
  assign n602 = pi043 & ~pi203;
  assign n603 = ~pi044 & pi204;
  assign n604 = pi044 & ~pi204;
  assign n605 = pi046 & ~pi206;
  assign n606 = pi045 & ~pi205;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~pi045 & pi205;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n604 & ~n609;
  assign n611 = ~n603 & ~n610;
  assign n612 = ~n602 & ~n611;
  assign n613 = ~n601 & ~n612;
  assign n614 = ~n600 & ~n613;
  assign n615 = ~n599 & ~n614;
  assign n616 = ~pi041 & ~n615;
  assign n617 = pi041 & ~n599;
  assign n618 = ~n614 & n617;
  assign n619 = pi201 & ~n618;
  assign n620 = ~pi040 & pi200;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n616 & n621;
  assign n623 = pi039 & ~pi199;
  assign n624 = pi040 & ~pi200;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n622 & n625;
  assign n627 = ~n598 & ~n626;
  assign n628 = ~pi039 & pi207;
  assign n629 = ~pi042 & pi210;
  assign n630 = pi042 & ~pi210;
  assign n631 = ~pi043 & pi211;
  assign n632 = pi043 & ~pi211;
  assign n633 = ~pi044 & pi212;
  assign n634 = pi044 & ~pi212;
  assign n635 = pi046 & ~pi214;
  assign n636 = pi045 & ~pi213;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~pi045 & pi213;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n634 & ~n639;
  assign n641 = ~n633 & ~n640;
  assign n642 = ~n632 & ~n641;
  assign n643 = ~n631 & ~n642;
  assign n644 = ~n630 & ~n643;
  assign n645 = ~n629 & ~n644;
  assign n646 = ~pi041 & ~n645;
  assign n647 = pi041 & ~n629;
  assign n648 = ~n644 & n647;
  assign n649 = pi209 & ~n648;
  assign n650 = ~pi040 & pi208;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n646 & n651;
  assign n653 = pi039 & ~pi207;
  assign n654 = pi040 & ~pi208;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n652 & n655;
  assign n657 = ~n628 & ~n656;
  assign n658 = ~n627 & ~n657;
  assign n659 = ~pi039 & pi239;
  assign n660 = ~pi042 & pi242;
  assign n661 = pi042 & ~pi242;
  assign n662 = ~pi043 & pi243;
  assign n663 = pi043 & ~pi243;
  assign n664 = ~pi044 & pi244;
  assign n665 = pi044 & ~pi244;
  assign n666 = pi046 & ~pi246;
  assign n667 = pi045 & ~pi245;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~pi045 & pi245;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~n665 & ~n670;
  assign n672 = ~n664 & ~n671;
  assign n673 = ~n663 & ~n672;
  assign n674 = ~n662 & ~n673;
  assign n675 = ~n661 & ~n674;
  assign n676 = ~n660 & ~n675;
  assign n677 = ~pi041 & ~n676;
  assign n678 = pi041 & ~n660;
  assign n679 = ~n675 & n678;
  assign n680 = pi241 & ~n679;
  assign n681 = ~pi040 & pi240;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~n677 & n682;
  assign n684 = pi039 & ~pi239;
  assign n685 = pi040 & ~pi240;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n683 & n686;
  assign n688 = ~n659 & ~n687;
  assign n689 = ~pi039 & pi231;
  assign n690 = ~pi042 & pi234;
  assign n691 = pi042 & ~pi234;
  assign n692 = ~pi043 & pi235;
  assign n693 = pi043 & ~pi235;
  assign n694 = ~pi044 & pi236;
  assign n695 = pi044 & ~pi236;
  assign n696 = pi046 & ~pi238;
  assign n697 = pi045 & ~pi237;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~pi045 & pi237;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~n695 & ~n700;
  assign n702 = ~n694 & ~n701;
  assign n703 = ~n693 & ~n702;
  assign n704 = ~n692 & ~n703;
  assign n705 = ~n691 & ~n704;
  assign n706 = ~n690 & ~n705;
  assign n707 = ~pi041 & ~n706;
  assign n708 = pi041 & ~n690;
  assign n709 = ~n705 & n708;
  assign n710 = pi233 & ~n709;
  assign n711 = ~pi040 & pi232;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~n707 & n712;
  assign n714 = pi040 & ~pi232;
  assign n715 = pi039 & ~pi231;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n713 & n716;
  assign n718 = ~n689 & ~n717;
  assign n719 = ~n688 & ~n718;
  assign n720 = n658 & n719;
  assign n721 = ~pi039 & pi247;
  assign n722 = ~pi042 & pi250;
  assign n723 = pi042 & ~pi250;
  assign n724 = ~pi043 & pi251;
  assign n725 = pi043 & ~pi251;
  assign n726 = ~pi044 & pi252;
  assign n727 = pi044 & ~pi252;
  assign n728 = pi046 & ~pi254;
  assign n729 = pi045 & ~pi253;
  assign n730 = ~n728 & ~n729;
  assign n731 = ~pi045 & pi253;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n727 & ~n732;
  assign n734 = ~n726 & ~n733;
  assign n735 = ~n725 & ~n734;
  assign n736 = ~n724 & ~n735;
  assign n737 = ~n723 & ~n736;
  assign n738 = ~n722 & ~n737;
  assign n739 = ~pi041 & ~n738;
  assign n740 = pi041 & ~n722;
  assign n741 = ~n737 & n740;
  assign n742 = pi249 & ~n741;
  assign n743 = ~pi040 & pi248;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n739 & n744;
  assign n746 = pi039 & ~pi247;
  assign n747 = pi040 & ~pi248;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n745 & n748;
  assign n750 = ~n721 & ~n749;
  assign n751 = ~pi039 & pi263;
  assign n752 = ~pi042 & pi266;
  assign n753 = pi042 & ~pi266;
  assign n754 = ~pi043 & pi267;
  assign n755 = pi043 & ~pi267;
  assign n756 = ~pi044 & pi268;
  assign n757 = pi044 & ~pi268;
  assign n758 = pi046 & ~pi270;
  assign n759 = pi045 & ~pi269;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~pi045 & pi269;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n757 & ~n762;
  assign n764 = ~n756 & ~n763;
  assign n765 = ~n755 & ~n764;
  assign n766 = ~n754 & ~n765;
  assign n767 = ~n753 & ~n766;
  assign n768 = ~n752 & ~n767;
  assign n769 = ~pi041 & ~n768;
  assign n770 = pi041 & ~n752;
  assign n771 = ~n767 & n770;
  assign n772 = pi265 & ~n771;
  assign n773 = ~pi040 & pi264;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n769 & n774;
  assign n776 = pi039 & ~pi263;
  assign n777 = pi040 & ~pi264;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n775 & n778;
  assign n780 = ~n751 & ~n779;
  assign n781 = ~n750 & ~n780;
  assign n782 = ~pi039 & pi223;
  assign n783 = ~pi042 & pi226;
  assign n784 = pi042 & ~pi226;
  assign n785 = ~pi043 & pi227;
  assign n786 = pi043 & ~pi227;
  assign n787 = ~pi044 & pi228;
  assign n788 = pi044 & ~pi228;
  assign n789 = pi046 & ~pi230;
  assign n790 = pi045 & ~pi229;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~pi045 & pi229;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n788 & ~n793;
  assign n795 = ~n787 & ~n794;
  assign n796 = ~n786 & ~n795;
  assign n797 = ~n785 & ~n796;
  assign n798 = ~n784 & ~n797;
  assign n799 = ~n783 & ~n798;
  assign n800 = ~pi041 & ~n799;
  assign n801 = pi041 & ~n783;
  assign n802 = ~n798 & n801;
  assign n803 = pi225 & ~n802;
  assign n804 = ~pi040 & pi224;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n800 & n805;
  assign n807 = pi039 & ~pi223;
  assign n808 = pi040 & ~pi224;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n806 & n809;
  assign n811 = ~n782 & ~n810;
  assign n812 = ~pi039 & pi215;
  assign n813 = ~pi042 & pi218;
  assign n814 = pi042 & ~pi218;
  assign n815 = ~pi043 & pi219;
  assign n816 = pi043 & ~pi219;
  assign n817 = ~pi044 & pi220;
  assign n818 = pi044 & ~pi220;
  assign n819 = pi046 & ~pi222;
  assign n820 = pi045 & ~pi221;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~pi045 & pi221;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n818 & ~n823;
  assign n825 = ~n817 & ~n824;
  assign n826 = ~n816 & ~n825;
  assign n827 = ~n815 & ~n826;
  assign n828 = ~n814 & ~n827;
  assign n829 = ~n813 & ~n828;
  assign n830 = ~pi041 & ~n829;
  assign n831 = pi041 & ~n813;
  assign n832 = ~n828 & n831;
  assign n833 = pi217 & ~n832;
  assign n834 = ~pi040 & pi216;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~n830 & n835;
  assign n837 = pi039 & ~pi215;
  assign n838 = pi040 & ~pi216;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n836 & n839;
  assign n841 = ~n812 & ~n840;
  assign n842 = ~n811 & ~n841;
  assign n843 = n781 & n842;
  assign n844 = n720 & n843;
  assign n845 = n597 & n844;
  assign n846 = ~pi039 & pi103;
  assign n847 = pi039 & ~pi103;
  assign n848 = ~pi040 & pi104;
  assign n849 = pi040 & ~pi104;
  assign n850 = pi042 & ~pi106;
  assign n851 = ~pi043 & pi107;
  assign n852 = pi043 & ~pi107;
  assign n853 = ~pi044 & pi108;
  assign n854 = pi044 & ~pi108;
  assign n855 = pi046 & ~pi110;
  assign n856 = pi045 & ~pi109;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~pi045 & pi109;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n854 & ~n859;
  assign n861 = ~n853 & ~n860;
  assign n862 = ~n852 & ~n861;
  assign n863 = ~n851 & ~n862;
  assign n864 = ~n850 & ~n863;
  assign n865 = ~pi042 & pi106;
  assign n866 = pi041 & ~n865;
  assign n867 = ~n864 & n866;
  assign n868 = pi105 & ~n867;
  assign n869 = ~n864 & ~n865;
  assign n870 = ~pi041 & ~n869;
  assign n871 = ~n868 & ~n870;
  assign n872 = ~n849 & ~n871;
  assign n873 = ~n848 & ~n872;
  assign n874 = ~n847 & ~n873;
  assign n875 = ~n846 & ~n874;
  assign n876 = ~pi039 & pi071;
  assign n877 = pi039 & ~pi071;
  assign n878 = ~pi040 & pi072;
  assign n879 = pi040 & ~pi072;
  assign n880 = pi042 & ~pi074;
  assign n881 = ~pi043 & pi075;
  assign n882 = pi043 & ~pi075;
  assign n883 = ~pi044 & pi076;
  assign n884 = pi044 & ~pi076;
  assign n885 = pi046 & ~pi078;
  assign n886 = pi045 & ~pi077;
  assign n887 = ~n885 & ~n886;
  assign n888 = ~pi045 & pi077;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n884 & ~n889;
  assign n891 = ~n883 & ~n890;
  assign n892 = ~n882 & ~n891;
  assign n893 = ~n881 & ~n892;
  assign n894 = ~n880 & ~n893;
  assign n895 = ~pi042 & pi074;
  assign n896 = pi041 & ~n895;
  assign n897 = ~n894 & n896;
  assign n898 = pi073 & ~n897;
  assign n899 = ~n894 & ~n895;
  assign n900 = ~pi041 & ~n899;
  assign n901 = ~n898 & ~n900;
  assign n902 = ~n879 & ~n901;
  assign n903 = ~n878 & ~n902;
  assign n904 = ~n877 & ~n903;
  assign n905 = ~n876 & ~n904;
  assign n906 = ~n875 & ~n905;
  assign n907 = ~pi039 & pi055;
  assign n908 = pi039 & ~pi055;
  assign n909 = ~pi040 & pi056;
  assign n910 = pi040 & ~pi056;
  assign n911 = pi042 & ~pi058;
  assign n912 = ~pi043 & pi059;
  assign n913 = pi043 & ~pi059;
  assign n914 = ~pi044 & pi060;
  assign n915 = pi044 & ~pi060;
  assign n916 = pi046 & ~pi062;
  assign n917 = pi045 & ~pi061;
  assign n918 = ~n916 & ~n917;
  assign n919 = ~pi045 & pi061;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n915 & ~n920;
  assign n922 = ~n914 & ~n921;
  assign n923 = ~n913 & ~n922;
  assign n924 = ~n912 & ~n923;
  assign n925 = ~n911 & ~n924;
  assign n926 = ~pi042 & pi058;
  assign n927 = pi041 & ~n926;
  assign n928 = ~n925 & n927;
  assign n929 = pi057 & ~n928;
  assign n930 = ~n925 & ~n926;
  assign n931 = ~pi041 & ~n930;
  assign n932 = ~n929 & ~n931;
  assign n933 = ~n910 & ~n932;
  assign n934 = ~n909 & ~n933;
  assign n935 = ~n908 & ~n934;
  assign n936 = ~n907 & ~n935;
  assign n937 = ~pi039 & pi087;
  assign n938 = pi039 & ~pi087;
  assign n939 = ~pi040 & pi088;
  assign n940 = pi040 & ~pi088;
  assign n941 = pi042 & ~pi090;
  assign n942 = ~pi043 & pi091;
  assign n943 = pi043 & ~pi091;
  assign n944 = ~pi044 & pi092;
  assign n945 = pi044 & ~pi092;
  assign n946 = pi046 & ~pi094;
  assign n947 = pi045 & ~pi093;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~pi045 & pi093;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n945 & ~n950;
  assign n952 = ~n944 & ~n951;
  assign n953 = ~n943 & ~n952;
  assign n954 = ~n942 & ~n953;
  assign n955 = ~n941 & ~n954;
  assign n956 = ~pi042 & pi090;
  assign n957 = pi041 & ~n956;
  assign n958 = ~n955 & n957;
  assign n959 = pi089 & ~n958;
  assign n960 = ~n955 & ~n956;
  assign n961 = ~pi041 & ~n960;
  assign n962 = ~n959 & ~n961;
  assign n963 = ~n940 & ~n962;
  assign n964 = ~n939 & ~n963;
  assign n965 = ~n938 & ~n964;
  assign n966 = ~n937 & ~n965;
  assign n967 = ~n936 & ~n966;
  assign n968 = n906 & n967;
  assign n969 = ~pi039 & pi111;
  assign n970 = pi043 & ~pi115;
  assign n971 = ~pi043 & pi115;
  assign n972 = pi045 & ~pi117;
  assign n973 = ~pi045 & pi117;
  assign n974 = pi046 & ~pi118;
  assign n975 = ~n973 & n974;
  assign n976 = ~n972 & ~n975;
  assign n977 = ~pi044 & pi116;
  assign n978 = ~n976 & ~n977;
  assign n979 = pi044 & ~pi116;
  assign n980 = ~n978 & ~n979;
  assign n981 = ~n971 & ~n980;
  assign n982 = ~n970 & ~n981;
  assign n983 = ~pi042 & pi114;
  assign n984 = ~n982 & ~n983;
  assign n985 = pi042 & ~pi114;
  assign n986 = pi041 & ~pi113;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n984 & n987;
  assign n989 = ~pi040 & pi112;
  assign n990 = ~pi041 & pi113;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n988 & n991;
  assign n993 = pi040 & ~pi112;
  assign n994 = pi039 & ~pi111;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~n992 & n995;
  assign n997 = ~n969 & ~n996;
  assign n998 = ~pi039 & pi167;
  assign n999 = pi043 & ~pi171;
  assign n1000 = ~pi043 & pi171;
  assign n1001 = pi045 & ~pi173;
  assign n1002 = ~pi045 & pi173;
  assign n1003 = pi046 & ~pi174;
  assign n1004 = ~n1002 & n1003;
  assign n1005 = ~n1001 & ~n1004;
  assign n1006 = ~pi044 & pi172;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = pi044 & ~pi172;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~n1000 & ~n1009;
  assign n1011 = ~n999 & ~n1010;
  assign n1012 = ~pi042 & pi170;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = pi042 & ~pi170;
  assign n1015 = pi041 & ~pi169;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n1013 & n1016;
  assign n1018 = ~pi040 & pi168;
  assign n1019 = ~pi041 & pi169;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~n1017 & n1020;
  assign n1022 = pi040 & ~pi168;
  assign n1023 = pi039 & ~pi167;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n1021 & n1024;
  assign n1026 = ~n998 & ~n1025;
  assign n1027 = ~pi039 & pi135;
  assign n1028 = pi043 & ~pi139;
  assign n1029 = ~pi043 & pi139;
  assign n1030 = pi045 & ~pi141;
  assign n1031 = ~pi045 & pi141;
  assign n1032 = pi046 & ~pi142;
  assign n1033 = ~n1031 & n1032;
  assign n1034 = ~n1030 & ~n1033;
  assign n1035 = ~pi044 & pi140;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = pi044 & ~pi140;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = ~n1029 & ~n1038;
  assign n1040 = ~n1028 & ~n1039;
  assign n1041 = ~pi042 & pi138;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = pi042 & ~pi138;
  assign n1044 = pi041 & ~pi137;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~n1042 & n1045;
  assign n1047 = ~pi040 & pi136;
  assign n1048 = ~pi041 & pi137;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = ~n1046 & n1049;
  assign n1051 = pi040 & ~pi136;
  assign n1052 = pi039 & ~pi135;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n1050 & n1053;
  assign n1055 = ~n1027 & ~n1054;
  assign n1056 = ~n1026 & ~n1055;
  assign n1057 = ~n997 & n1056;
  assign n1058 = ~pi039 & pi175;
  assign n1059 = pi039 & ~pi175;
  assign n1060 = ~pi040 & pi176;
  assign n1061 = pi040 & ~pi176;
  assign n1062 = ~pi041 & pi177;
  assign n1063 = pi043 & ~pi179;
  assign n1064 = ~pi043 & pi179;
  assign n1065 = pi044 & ~pi180;
  assign n1066 = pi045 & ~pi181;
  assign n1067 = pi046 & ~pi182;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~pi045 & pi181;
  assign n1070 = ~pi044 & pi180;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1068 & n1071;
  assign n1073 = ~n1065 & ~n1072;
  assign n1074 = ~n1064 & ~n1073;
  assign n1075 = ~n1063 & ~n1074;
  assign n1076 = ~pi042 & pi178;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = pi042 & ~pi178;
  assign n1079 = pi041 & ~pi177;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~n1077 & n1080;
  assign n1082 = ~n1062 & ~n1081;
  assign n1083 = ~n1061 & ~n1082;
  assign n1084 = ~n1060 & ~n1083;
  assign n1085 = ~n1059 & ~n1084;
  assign n1086 = ~n1058 & ~n1085;
  assign n1087 = ~pi039 & pi183;
  assign n1088 = pi043 & ~pi187;
  assign n1089 = ~pi043 & pi187;
  assign n1090 = pi045 & ~pi189;
  assign n1091 = ~pi045 & pi189;
  assign n1092 = pi046 & ~pi190;
  assign n1093 = ~n1091 & n1092;
  assign n1094 = ~n1090 & ~n1093;
  assign n1095 = ~pi044 & pi188;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = pi044 & ~pi188;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1089 & ~n1098;
  assign n1100 = ~n1088 & ~n1099;
  assign n1101 = ~pi042 & pi186;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = pi042 & ~pi186;
  assign n1104 = pi041 & ~pi185;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~n1102 & n1105;
  assign n1107 = ~pi040 & pi184;
  assign n1108 = ~pi041 & pi185;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~n1106 & n1109;
  assign n1111 = pi040 & ~pi184;
  assign n1112 = pi039 & ~pi183;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1110 & n1113;
  assign n1115 = ~n1087 & ~n1114;
  assign n1116 = ~pi039 & pi151;
  assign n1117 = pi043 & ~pi155;
  assign n1118 = ~pi043 & pi155;
  assign n1119 = pi044 & ~pi156;
  assign n1120 = pi045 & ~pi157;
  assign n1121 = pi046 & ~pi158;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~pi045 & pi157;
  assign n1124 = ~pi044 & pi156;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1122 & n1125;
  assign n1127 = ~n1119 & ~n1126;
  assign n1128 = ~n1118 & ~n1127;
  assign n1129 = ~n1117 & ~n1128;
  assign n1130 = ~pi042 & pi154;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = pi042 & ~pi154;
  assign n1133 = pi041 & ~pi153;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1131 & n1134;
  assign n1136 = ~pi040 & pi152;
  assign n1137 = ~pi041 & pi153;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = ~n1135 & n1138;
  assign n1140 = pi040 & ~pi152;
  assign n1141 = pi039 & ~pi151;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = ~n1139 & n1142;
  assign n1144 = ~n1116 & ~n1143;
  assign n1145 = ~pi039 & pi127;
  assign n1146 = pi043 & ~pi131;
  assign n1147 = ~pi045 & pi133;
  assign n1148 = pi046 & ~pi134;
  assign n1149 = ~n1147 & n1148;
  assign n1150 = pi045 & ~pi133;
  assign n1151 = pi044 & ~pi132;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n1149 & n1152;
  assign n1154 = ~pi044 & pi132;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = ~n1146 & ~n1155;
  assign n1157 = ~pi043 & pi131;
  assign n1158 = ~pi042 & pi130;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n1156 & n1159;
  assign n1161 = pi041 & ~pi129;
  assign n1162 = pi042 & ~pi130;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1160 & n1163;
  assign n1165 = ~pi040 & pi128;
  assign n1166 = ~pi041 & pi129;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1164 & n1167;
  assign n1169 = pi040 & ~pi128;
  assign n1170 = pi039 & ~pi127;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n1168 & n1171;
  assign n1173 = ~n1145 & ~n1172;
  assign n1174 = pi001 & ~n1173;
  assign n1175 = ~n1144 & n1174;
  assign n1176 = ~n1115 & n1175;
  assign n1177 = ~n1086 & n1176;
  assign n1178 = n1057 & n1177;
  assign n1179 = ~pi039 & pi271;
  assign n1180 = ~pi042 & pi274;
  assign n1181 = pi042 & ~pi274;
  assign n1182 = ~pi043 & pi275;
  assign n1183 = pi043 & ~pi275;
  assign n1184 = ~pi044 & pi276;
  assign n1185 = pi044 & ~pi276;
  assign n1186 = pi046 & ~pi278;
  assign n1187 = pi045 & ~pi277;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~pi045 & pi277;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = ~n1185 & ~n1190;
  assign n1192 = ~n1184 & ~n1191;
  assign n1193 = ~n1183 & ~n1192;
  assign n1194 = ~n1182 & ~n1193;
  assign n1195 = ~n1181 & ~n1194;
  assign n1196 = ~n1180 & ~n1195;
  assign n1197 = ~pi041 & ~n1196;
  assign n1198 = pi041 & ~n1180;
  assign n1199 = ~n1195 & n1198;
  assign n1200 = pi273 & ~n1199;
  assign n1201 = ~pi040 & pi272;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1197 & n1202;
  assign n1204 = pi039 & ~pi271;
  assign n1205 = pi040 & ~pi272;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n1203 & n1206;
  assign n1208 = ~n1179 & ~n1207;
  assign n1209 = ~pi039 & pi255;
  assign n1210 = ~pi042 & pi258;
  assign n1211 = pi042 & ~pi258;
  assign n1212 = ~pi043 & pi259;
  assign n1213 = pi043 & ~pi259;
  assign n1214 = ~pi044 & pi260;
  assign n1215 = pi044 & ~pi260;
  assign n1216 = pi046 & ~pi262;
  assign n1217 = pi045 & ~pi261;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~pi045 & pi261;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~n1215 & ~n1220;
  assign n1222 = ~n1214 & ~n1221;
  assign n1223 = ~n1213 & ~n1222;
  assign n1224 = ~n1212 & ~n1223;
  assign n1225 = ~n1211 & ~n1224;
  assign n1226 = ~n1210 & ~n1225;
  assign n1227 = ~pi041 & ~n1226;
  assign n1228 = pi041 & ~n1210;
  assign n1229 = ~n1225 & n1228;
  assign n1230 = pi257 & ~n1229;
  assign n1231 = ~pi040 & pi256;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1227 & n1232;
  assign n1234 = pi040 & ~pi256;
  assign n1235 = pi039 & ~pi255;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~n1233 & n1236;
  assign n1238 = ~n1209 & ~n1237;
  assign n1239 = ~n1208 & ~n1238;
  assign n1240 = n1178 & n1239;
  assign n1241 = ~pi039 & pi191;
  assign n1242 = pi039 & ~pi191;
  assign n1243 = ~pi040 & pi192;
  assign n1244 = pi040 & ~pi192;
  assign n1245 = pi042 & ~pi194;
  assign n1246 = ~pi043 & pi195;
  assign n1247 = pi043 & ~pi195;
  assign n1248 = ~pi044 & pi196;
  assign n1249 = pi044 & ~pi196;
  assign n1250 = pi046 & ~pi198;
  assign n1251 = pi045 & ~pi197;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~pi045 & pi197;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1249 & ~n1254;
  assign n1256 = ~n1248 & ~n1255;
  assign n1257 = ~n1247 & ~n1256;
  assign n1258 = ~n1246 & ~n1257;
  assign n1259 = ~n1245 & ~n1258;
  assign n1260 = ~pi042 & pi194;
  assign n1261 = pi041 & ~n1260;
  assign n1262 = ~n1259 & n1261;
  assign n1263 = pi193 & ~n1262;
  assign n1264 = ~n1259 & ~n1260;
  assign n1265 = ~pi041 & ~n1264;
  assign n1266 = ~n1263 & ~n1265;
  assign n1267 = ~n1244 & ~n1266;
  assign n1268 = ~n1243 & ~n1267;
  assign n1269 = ~n1242 & ~n1268;
  assign n1270 = ~n1241 & ~n1269;
  assign n1271 = ~pi039 & pi159;
  assign n1272 = pi039 & ~pi159;
  assign n1273 = ~pi040 & pi160;
  assign n1274 = pi040 & ~pi160;
  assign n1275 = ~pi041 & pi161;
  assign n1276 = pi043 & ~pi163;
  assign n1277 = ~pi043 & pi163;
  assign n1278 = pi044 & ~pi164;
  assign n1279 = pi045 & ~pi165;
  assign n1280 = pi046 & ~pi166;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~pi045 & pi165;
  assign n1283 = ~pi044 & pi164;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = ~n1281 & n1284;
  assign n1286 = ~n1278 & ~n1285;
  assign n1287 = ~n1277 & ~n1286;
  assign n1288 = ~n1276 & ~n1287;
  assign n1289 = ~pi042 & pi162;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = pi042 & ~pi162;
  assign n1292 = pi041 & ~pi161;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1290 & n1293;
  assign n1295 = ~n1275 & ~n1294;
  assign n1296 = ~n1274 & ~n1295;
  assign n1297 = ~n1273 & ~n1296;
  assign n1298 = ~n1272 & ~n1297;
  assign n1299 = ~n1271 & ~n1298;
  assign n1300 = ~pi039 & pi119;
  assign n1301 = pi039 & ~pi119;
  assign n1302 = ~pi040 & pi120;
  assign n1303 = pi040 & ~pi120;
  assign n1304 = ~pi041 & pi121;
  assign n1305 = pi043 & ~pi123;
  assign n1306 = ~pi043 & pi123;
  assign n1307 = pi044 & ~pi124;
  assign n1308 = pi045 & ~pi125;
  assign n1309 = pi046 & ~pi126;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~pi045 & pi125;
  assign n1312 = ~pi044 & pi124;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1310 & n1313;
  assign n1315 = ~n1307 & ~n1314;
  assign n1316 = ~n1306 & ~n1315;
  assign n1317 = ~n1305 & ~n1316;
  assign n1318 = ~pi042 & pi122;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = pi042 & ~pi122;
  assign n1321 = pi041 & ~pi121;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1319 & n1322;
  assign n1324 = ~n1304 & ~n1323;
  assign n1325 = ~n1303 & ~n1324;
  assign n1326 = ~n1302 & ~n1325;
  assign n1327 = ~n1301 & ~n1326;
  assign n1328 = ~n1300 & ~n1327;
  assign n1329 = ~pi039 & pi143;
  assign n1330 = pi039 & ~pi143;
  assign n1331 = ~pi040 & pi144;
  assign n1332 = pi040 & ~pi144;
  assign n1333 = ~pi041 & pi145;
  assign n1334 = pi043 & ~pi147;
  assign n1335 = ~pi043 & pi147;
  assign n1336 = pi044 & ~pi148;
  assign n1337 = pi045 & ~pi149;
  assign n1338 = pi046 & ~pi150;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~pi045 & pi149;
  assign n1341 = ~pi044 & pi148;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = ~n1339 & n1342;
  assign n1344 = ~n1336 & ~n1343;
  assign n1345 = ~n1335 & ~n1344;
  assign n1346 = ~n1334 & ~n1345;
  assign n1347 = ~pi042 & pi146;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = pi042 & ~pi146;
  assign n1350 = pi041 & ~pi145;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1348 & n1351;
  assign n1353 = ~n1333 & ~n1352;
  assign n1354 = ~n1332 & ~n1353;
  assign n1355 = ~n1331 & ~n1354;
  assign n1356 = ~n1330 & ~n1355;
  assign n1357 = ~n1329 & ~n1356;
  assign n1358 = ~n1328 & ~n1357;
  assign n1359 = ~n1299 & n1358;
  assign n1360 = ~n1270 & n1359;
  assign n1361 = n1240 & n1360;
  assign n1362 = n968 & n1361;
  assign n1363 = n845 & n1362;
  assign po001 = n503 | n1363;
  assign n1365 = ~n1144 & ~n1173;
  assign n1366 = ~n1115 & n1365;
  assign n1367 = ~n1086 & n1366;
  assign n1368 = n1057 & n1367;
  assign n1369 = n1239 & n1368;
  assign n1370 = n1360 & n1369;
  assign n1371 = n968 & n1370;
  assign n1372 = n845 & n1371;
  assign n1373 = ~n936 & ~n1372;
  assign n1374 = ~pi055 & pi151;
  assign n1375 = ~pi058 & pi154;
  assign n1376 = pi058 & ~pi154;
  assign n1377 = ~pi059 & pi155;
  assign n1378 = pi059 & ~pi155;
  assign n1379 = ~pi060 & pi156;
  assign n1380 = pi060 & ~pi156;
  assign n1381 = pi062 & ~pi158;
  assign n1382 = pi061 & ~pi157;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~pi061 & pi157;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n1380 & ~n1385;
  assign n1387 = ~n1379 & ~n1386;
  assign n1388 = ~n1378 & ~n1387;
  assign n1389 = ~n1377 & ~n1388;
  assign n1390 = ~n1376 & ~n1389;
  assign n1391 = ~n1375 & ~n1390;
  assign n1392 = pi153 & ~n1391;
  assign n1393 = ~pi153 & ~n1375;
  assign n1394 = ~n1390 & n1393;
  assign n1395 = ~pi057 & ~n1394;
  assign n1396 = ~pi056 & pi152;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1392 & n1397;
  assign n1399 = pi056 & ~pi152;
  assign n1400 = pi055 & ~pi151;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1398 & n1401;
  assign n1403 = ~n1374 & ~n1402;
  assign n1404 = ~pi055 & pi111;
  assign n1405 = ~pi058 & pi114;
  assign n1406 = pi058 & ~pi114;
  assign n1407 = ~pi059 & pi115;
  assign n1408 = pi059 & ~pi115;
  assign n1409 = ~pi060 & pi116;
  assign n1410 = pi060 & ~pi116;
  assign n1411 = pi062 & ~pi118;
  assign n1412 = pi061 & ~pi117;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = ~pi061 & pi117;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~n1410 & ~n1415;
  assign n1417 = ~n1409 & ~n1416;
  assign n1418 = ~n1408 & ~n1417;
  assign n1419 = ~n1407 & ~n1418;
  assign n1420 = ~n1406 & ~n1419;
  assign n1421 = ~n1405 & ~n1420;
  assign n1422 = pi113 & ~n1421;
  assign n1423 = ~pi113 & ~n1405;
  assign n1424 = ~n1420 & n1423;
  assign n1425 = ~pi057 & ~n1424;
  assign n1426 = ~pi056 & pi112;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1422 & n1427;
  assign n1429 = pi056 & ~pi112;
  assign n1430 = pi055 & ~pi111;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1428 & n1431;
  assign n1433 = ~n1404 & ~n1432;
  assign n1434 = ~n1403 & ~n1433;
  assign n1435 = ~pi055 & pi079;
  assign n1436 = ~pi058 & pi082;
  assign n1437 = pi058 & ~pi082;
  assign n1438 = ~pi059 & pi083;
  assign n1439 = pi059 & ~pi083;
  assign n1440 = ~pi060 & pi084;
  assign n1441 = pi060 & ~pi084;
  assign n1442 = pi062 & ~pi086;
  assign n1443 = pi061 & ~pi085;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~pi061 & pi085;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = ~n1441 & ~n1446;
  assign n1448 = ~n1440 & ~n1447;
  assign n1449 = ~n1439 & ~n1448;
  assign n1450 = ~n1438 & ~n1449;
  assign n1451 = ~n1437 & ~n1450;
  assign n1452 = ~n1436 & ~n1451;
  assign n1453 = ~pi057 & ~n1452;
  assign n1454 = pi057 & ~n1436;
  assign n1455 = ~n1451 & n1454;
  assign n1456 = pi081 & ~n1455;
  assign n1457 = ~pi056 & pi080;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1453 & n1458;
  assign n1460 = pi056 & ~pi080;
  assign n1461 = pi055 & ~pi079;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~n1459 & n1462;
  assign n1464 = ~n1435 & ~n1463;
  assign n1465 = ~pi055 & pi063;
  assign n1466 = ~pi058 & pi066;
  assign n1467 = pi058 & ~pi066;
  assign n1468 = ~pi059 & pi067;
  assign n1469 = pi059 & ~pi067;
  assign n1470 = ~pi060 & pi068;
  assign n1471 = pi060 & ~pi068;
  assign n1472 = pi062 & ~pi070;
  assign n1473 = pi061 & ~pi069;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = ~pi061 & pi069;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~n1471 & ~n1476;
  assign n1478 = ~n1470 & ~n1477;
  assign n1479 = ~n1469 & ~n1478;
  assign n1480 = ~n1468 & ~n1479;
  assign n1481 = ~n1467 & ~n1480;
  assign n1482 = ~n1466 & ~n1481;
  assign n1483 = ~pi057 & ~n1482;
  assign n1484 = pi057 & ~n1466;
  assign n1485 = ~n1481 & n1484;
  assign n1486 = pi065 & ~n1485;
  assign n1487 = ~pi056 & pi064;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1483 & n1488;
  assign n1490 = pi056 & ~pi064;
  assign n1491 = pi055 & ~pi063;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1489 & n1492;
  assign n1494 = ~n1465 & ~n1493;
  assign n1495 = ~n1464 & ~n1494;
  assign n1496 = n1434 & n1495;
  assign n1497 = ~pi055 & pi271;
  assign n1498 = ~pi058 & pi274;
  assign n1499 = pi058 & ~pi274;
  assign n1500 = ~pi059 & pi275;
  assign n1501 = pi059 & ~pi275;
  assign n1502 = ~pi060 & pi276;
  assign n1503 = pi060 & ~pi276;
  assign n1504 = pi062 & ~pi278;
  assign n1505 = pi061 & ~pi277;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = ~pi061 & pi277;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1503 & ~n1508;
  assign n1510 = ~n1502 & ~n1509;
  assign n1511 = ~n1501 & ~n1510;
  assign n1512 = ~n1500 & ~n1511;
  assign n1513 = ~n1499 & ~n1512;
  assign n1514 = ~n1498 & ~n1513;
  assign n1515 = pi273 & ~n1514;
  assign n1516 = ~pi273 & ~n1498;
  assign n1517 = ~n1513 & n1516;
  assign n1518 = ~pi057 & ~n1517;
  assign n1519 = ~pi056 & pi272;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = ~n1515 & n1520;
  assign n1522 = pi056 & ~pi272;
  assign n1523 = pi055 & ~pi271;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1521 & n1524;
  assign n1526 = ~n1497 & ~n1525;
  assign n1527 = ~pi055 & pi263;
  assign n1528 = ~pi058 & pi266;
  assign n1529 = pi058 & ~pi266;
  assign n1530 = ~pi059 & pi267;
  assign n1531 = pi059 & ~pi267;
  assign n1532 = ~pi060 & pi268;
  assign n1533 = pi060 & ~pi268;
  assign n1534 = pi062 & ~pi270;
  assign n1535 = pi061 & ~pi269;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~pi061 & pi269;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1533 & ~n1538;
  assign n1540 = ~n1532 & ~n1539;
  assign n1541 = ~n1531 & ~n1540;
  assign n1542 = ~n1530 & ~n1541;
  assign n1543 = ~n1529 & ~n1542;
  assign n1544 = ~n1528 & ~n1543;
  assign n1545 = pi265 & ~n1544;
  assign n1546 = ~pi265 & ~n1528;
  assign n1547 = ~n1543 & n1546;
  assign n1548 = ~pi057 & ~n1547;
  assign n1549 = ~pi056 & pi264;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~n1545 & n1550;
  assign n1552 = pi056 & ~pi264;
  assign n1553 = pi055 & ~pi263;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1551 & n1554;
  assign n1556 = ~n1527 & ~n1555;
  assign n1557 = ~n1526 & ~n1556;
  assign n1558 = ~pi055 & pi247;
  assign n1559 = ~pi058 & pi250;
  assign n1560 = pi058 & ~pi250;
  assign n1561 = ~pi059 & pi251;
  assign n1562 = pi059 & ~pi251;
  assign n1563 = ~pi060 & pi252;
  assign n1564 = pi060 & ~pi252;
  assign n1565 = pi062 & ~pi254;
  assign n1566 = pi061 & ~pi253;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~pi061 & pi253;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = ~n1564 & ~n1569;
  assign n1571 = ~n1563 & ~n1570;
  assign n1572 = ~n1562 & ~n1571;
  assign n1573 = ~n1561 & ~n1572;
  assign n1574 = ~n1560 & ~n1573;
  assign n1575 = ~n1559 & ~n1574;
  assign n1576 = pi249 & ~n1575;
  assign n1577 = ~pi249 & ~n1559;
  assign n1578 = ~n1574 & n1577;
  assign n1579 = ~pi057 & ~n1578;
  assign n1580 = ~pi056 & pi248;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1576 & n1581;
  assign n1583 = pi056 & ~pi248;
  assign n1584 = pi055 & ~pi247;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = ~n1582 & n1585;
  assign n1587 = ~n1558 & ~n1586;
  assign n1588 = ~pi055 & pi215;
  assign n1589 = ~pi058 & pi218;
  assign n1590 = pi058 & ~pi218;
  assign n1591 = ~pi059 & pi219;
  assign n1592 = pi059 & ~pi219;
  assign n1593 = ~pi060 & pi220;
  assign n1594 = pi060 & ~pi220;
  assign n1595 = pi062 & ~pi222;
  assign n1596 = pi061 & ~pi221;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~pi061 & pi221;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1594 & ~n1599;
  assign n1601 = ~n1593 & ~n1600;
  assign n1602 = ~n1592 & ~n1601;
  assign n1603 = ~n1591 & ~n1602;
  assign n1604 = ~n1590 & ~n1603;
  assign n1605 = ~n1589 & ~n1604;
  assign n1606 = pi217 & ~n1605;
  assign n1607 = ~pi217 & ~n1589;
  assign n1608 = ~n1604 & n1607;
  assign n1609 = ~pi057 & ~n1608;
  assign n1610 = ~pi056 & pi216;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1606 & n1611;
  assign n1613 = pi056 & ~pi216;
  assign n1614 = pi055 & ~pi215;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = ~n1588 & ~n1616;
  assign n1618 = ~n1587 & ~n1617;
  assign n1619 = n1557 & n1618;
  assign n1620 = ~pi055 & pi183;
  assign n1621 = ~pi058 & pi186;
  assign n1622 = pi058 & ~pi186;
  assign n1623 = ~pi059 & pi187;
  assign n1624 = pi059 & ~pi187;
  assign n1625 = ~pi060 & pi188;
  assign n1626 = pi060 & ~pi188;
  assign n1627 = pi062 & ~pi190;
  assign n1628 = pi061 & ~pi189;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~pi061 & pi189;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n1626 & ~n1631;
  assign n1633 = ~n1625 & ~n1632;
  assign n1634 = ~n1624 & ~n1633;
  assign n1635 = ~n1623 & ~n1634;
  assign n1636 = ~n1622 & ~n1635;
  assign n1637 = ~n1621 & ~n1636;
  assign n1638 = pi185 & ~n1637;
  assign n1639 = ~pi185 & ~n1621;
  assign n1640 = ~n1636 & n1639;
  assign n1641 = ~pi057 & ~n1640;
  assign n1642 = ~pi056 & pi184;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1638 & n1643;
  assign n1645 = pi056 & ~pi184;
  assign n1646 = pi055 & ~pi183;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n1644 & n1647;
  assign n1649 = ~n1620 & ~n1648;
  assign n1650 = ~pi055 & pi239;
  assign n1651 = ~pi058 & pi242;
  assign n1652 = pi058 & ~pi242;
  assign n1653 = ~pi059 & pi243;
  assign n1654 = pi059 & ~pi243;
  assign n1655 = ~pi060 & pi244;
  assign n1656 = pi060 & ~pi244;
  assign n1657 = pi062 & ~pi246;
  assign n1658 = pi061 & ~pi245;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = ~pi061 & pi245;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~n1656 & ~n1661;
  assign n1663 = ~n1655 & ~n1662;
  assign n1664 = ~n1654 & ~n1663;
  assign n1665 = ~n1653 & ~n1664;
  assign n1666 = ~n1652 & ~n1665;
  assign n1667 = ~n1651 & ~n1666;
  assign n1668 = pi241 & ~n1667;
  assign n1669 = ~pi241 & ~n1651;
  assign n1670 = ~n1666 & n1669;
  assign n1671 = ~pi057 & ~n1670;
  assign n1672 = ~pi056 & pi240;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~n1668 & n1673;
  assign n1675 = pi056 & ~pi240;
  assign n1676 = pi055 & ~pi239;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = ~n1674 & n1677;
  assign n1679 = ~n1650 & ~n1678;
  assign n1680 = ~n1649 & ~n1679;
  assign n1681 = ~pi055 & pi231;
  assign n1682 = ~pi058 & pi234;
  assign n1683 = pi058 & ~pi234;
  assign n1684 = ~pi059 & pi235;
  assign n1685 = pi059 & ~pi235;
  assign n1686 = ~pi060 & pi236;
  assign n1687 = pi060 & ~pi236;
  assign n1688 = pi062 & ~pi238;
  assign n1689 = pi061 & ~pi237;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = ~pi061 & pi237;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1687 & ~n1692;
  assign n1694 = ~n1686 & ~n1693;
  assign n1695 = ~n1685 & ~n1694;
  assign n1696 = ~n1684 & ~n1695;
  assign n1697 = ~n1683 & ~n1696;
  assign n1698 = ~n1682 & ~n1697;
  assign n1699 = pi233 & ~n1698;
  assign n1700 = ~pi233 & ~n1682;
  assign n1701 = ~n1697 & n1700;
  assign n1702 = ~pi057 & ~n1701;
  assign n1703 = ~pi056 & pi232;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = ~n1699 & n1704;
  assign n1706 = pi056 & ~pi232;
  assign n1707 = pi055 & ~pi231;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n1705 & n1708;
  assign n1710 = ~n1681 & ~n1709;
  assign n1711 = ~pi055 & pi255;
  assign n1712 = ~pi058 & pi258;
  assign n1713 = pi058 & ~pi258;
  assign n1714 = ~pi059 & pi259;
  assign n1715 = pi059 & ~pi259;
  assign n1716 = ~pi060 & pi260;
  assign n1717 = pi060 & ~pi260;
  assign n1718 = pi062 & ~pi262;
  assign n1719 = pi061 & ~pi261;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~pi061 & pi261;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = ~n1717 & ~n1722;
  assign n1724 = ~n1716 & ~n1723;
  assign n1725 = ~n1715 & ~n1724;
  assign n1726 = ~n1714 & ~n1725;
  assign n1727 = ~n1713 & ~n1726;
  assign n1728 = ~n1712 & ~n1727;
  assign n1729 = pi257 & ~n1728;
  assign n1730 = ~pi257 & ~n1712;
  assign n1731 = ~n1727 & n1730;
  assign n1732 = ~pi057 & ~n1731;
  assign n1733 = ~pi056 & pi256;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~n1729 & n1734;
  assign n1736 = pi056 & ~pi256;
  assign n1737 = pi055 & ~pi255;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = ~n1711 & ~n1739;
  assign n1741 = ~n1710 & ~n1740;
  assign n1742 = n1680 & n1741;
  assign n1743 = n1619 & n1742;
  assign n1744 = n1496 & n1743;
  assign n1745 = ~pi055 & pi071;
  assign n1746 = pi055 & ~pi071;
  assign n1747 = ~pi056 & pi072;
  assign n1748 = pi056 & ~pi072;
  assign n1749 = pi058 & ~pi074;
  assign n1750 = ~pi059 & pi075;
  assign n1751 = pi059 & ~pi075;
  assign n1752 = ~pi060 & pi076;
  assign n1753 = pi060 & ~pi076;
  assign n1754 = pi062 & ~pi078;
  assign n1755 = pi061 & ~pi077;
  assign n1756 = ~n1754 & ~n1755;
  assign n1757 = ~pi061 & pi077;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~n1753 & ~n1758;
  assign n1760 = ~n1752 & ~n1759;
  assign n1761 = ~n1751 & ~n1760;
  assign n1762 = ~n1750 & ~n1761;
  assign n1763 = ~n1749 & ~n1762;
  assign n1764 = ~pi058 & pi074;
  assign n1765 = pi057 & ~n1764;
  assign n1766 = ~n1763 & n1765;
  assign n1767 = pi073 & ~n1766;
  assign n1768 = ~n1763 & ~n1764;
  assign n1769 = ~pi057 & ~n1768;
  assign n1770 = ~n1767 & ~n1769;
  assign n1771 = ~n1748 & ~n1770;
  assign n1772 = ~n1747 & ~n1771;
  assign n1773 = ~n1746 & ~n1772;
  assign n1774 = ~n1745 & ~n1773;
  assign n1775 = ~pi055 & pi159;
  assign n1776 = pi055 & ~pi159;
  assign n1777 = ~pi056 & pi160;
  assign n1778 = pi056 & ~pi160;
  assign n1779 = pi058 & ~pi162;
  assign n1780 = ~pi059 & pi163;
  assign n1781 = pi059 & ~pi163;
  assign n1782 = ~pi060 & pi164;
  assign n1783 = pi060 & ~pi164;
  assign n1784 = pi062 & ~pi166;
  assign n1785 = pi061 & ~pi165;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~pi061 & pi165;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = ~n1783 & ~n1788;
  assign n1790 = ~n1782 & ~n1789;
  assign n1791 = ~n1781 & ~n1790;
  assign n1792 = ~n1780 & ~n1791;
  assign n1793 = ~n1779 & ~n1792;
  assign n1794 = ~pi058 & pi162;
  assign n1795 = ~pi161 & ~n1794;
  assign n1796 = ~n1793 & n1795;
  assign n1797 = ~pi057 & ~n1796;
  assign n1798 = ~n1793 & ~n1794;
  assign n1799 = pi161 & ~n1798;
  assign n1800 = ~n1797 & ~n1799;
  assign n1801 = ~n1778 & ~n1800;
  assign n1802 = ~n1777 & ~n1801;
  assign n1803 = ~n1776 & ~n1802;
  assign n1804 = ~n1775 & ~n1803;
  assign n1805 = ~n1774 & ~n1804;
  assign n1806 = ~pi055 & pi103;
  assign n1807 = pi055 & ~pi103;
  assign n1808 = ~pi056 & pi104;
  assign n1809 = pi056 & ~pi104;
  assign n1810 = pi058 & ~pi106;
  assign n1811 = ~pi059 & pi107;
  assign n1812 = pi059 & ~pi107;
  assign n1813 = ~pi060 & pi108;
  assign n1814 = pi060 & ~pi108;
  assign n1815 = pi062 & ~pi110;
  assign n1816 = pi061 & ~pi109;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~pi061 & pi109;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~n1814 & ~n1819;
  assign n1821 = ~n1813 & ~n1820;
  assign n1822 = ~n1812 & ~n1821;
  assign n1823 = ~n1811 & ~n1822;
  assign n1824 = ~n1810 & ~n1823;
  assign n1825 = ~pi058 & pi106;
  assign n1826 = pi057 & ~n1825;
  assign n1827 = ~n1824 & n1826;
  assign n1828 = pi105 & ~n1827;
  assign n1829 = ~n1824 & ~n1825;
  assign n1830 = ~pi057 & ~n1829;
  assign n1831 = ~n1828 & ~n1830;
  assign n1832 = ~n1809 & ~n1831;
  assign n1833 = ~n1808 & ~n1832;
  assign n1834 = ~n1807 & ~n1833;
  assign n1835 = ~n1806 & ~n1834;
  assign n1836 = ~pi055 & pi087;
  assign n1837 = pi055 & ~pi087;
  assign n1838 = ~pi056 & pi088;
  assign n1839 = pi056 & ~pi088;
  assign n1840 = pi058 & ~pi090;
  assign n1841 = ~pi059 & pi091;
  assign n1842 = pi059 & ~pi091;
  assign n1843 = ~pi060 & pi092;
  assign n1844 = pi060 & ~pi092;
  assign n1845 = pi062 & ~pi094;
  assign n1846 = pi061 & ~pi093;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = ~pi061 & pi093;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1844 & ~n1849;
  assign n1851 = ~n1843 & ~n1850;
  assign n1852 = ~n1842 & ~n1851;
  assign n1853 = ~n1841 & ~n1852;
  assign n1854 = ~n1840 & ~n1853;
  assign n1855 = ~pi058 & pi090;
  assign n1856 = pi057 & ~n1855;
  assign n1857 = ~n1854 & n1856;
  assign n1858 = pi089 & ~n1857;
  assign n1859 = ~n1854 & ~n1855;
  assign n1860 = ~pi057 & ~n1859;
  assign n1861 = ~n1858 & ~n1860;
  assign n1862 = ~n1839 & ~n1861;
  assign n1863 = ~n1838 & ~n1862;
  assign n1864 = ~n1837 & ~n1863;
  assign n1865 = ~n1836 & ~n1864;
  assign n1866 = ~n1835 & ~n1865;
  assign n1867 = n1805 & n1866;
  assign n1868 = ~pi055 & pi191;
  assign n1869 = pi055 & ~pi191;
  assign n1870 = ~pi056 & pi192;
  assign n1871 = pi056 & ~pi192;
  assign n1872 = pi058 & ~pi194;
  assign n1873 = ~pi059 & pi195;
  assign n1874 = pi059 & ~pi195;
  assign n1875 = ~pi060 & pi196;
  assign n1876 = pi060 & ~pi196;
  assign n1877 = pi062 & ~pi198;
  assign n1878 = pi061 & ~pi197;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = ~pi061 & pi197;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~n1876 & ~n1881;
  assign n1883 = ~n1875 & ~n1882;
  assign n1884 = ~n1874 & ~n1883;
  assign n1885 = ~n1873 & ~n1884;
  assign n1886 = ~n1872 & ~n1885;
  assign n1887 = ~pi058 & pi194;
  assign n1888 = ~pi193 & ~n1887;
  assign n1889 = ~n1886 & n1888;
  assign n1890 = ~pi057 & ~n1889;
  assign n1891 = ~n1886 & ~n1887;
  assign n1892 = pi193 & ~n1891;
  assign n1893 = ~n1890 & ~n1892;
  assign n1894 = ~n1871 & ~n1893;
  assign n1895 = ~n1870 & ~n1894;
  assign n1896 = ~n1869 & ~n1895;
  assign n1897 = ~n1868 & ~n1896;
  assign n1898 = ~pi055 & pi143;
  assign n1899 = pi055 & ~pi143;
  assign n1900 = ~pi056 & pi144;
  assign n1901 = pi056 & ~pi144;
  assign n1902 = pi058 & ~pi146;
  assign n1903 = ~pi059 & pi147;
  assign n1904 = pi059 & ~pi147;
  assign n1905 = ~pi060 & pi148;
  assign n1906 = pi060 & ~pi148;
  assign n1907 = pi062 & ~pi150;
  assign n1908 = pi061 & ~pi149;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = ~pi061 & pi149;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1906 & ~n1911;
  assign n1913 = ~n1905 & ~n1912;
  assign n1914 = ~n1904 & ~n1913;
  assign n1915 = ~n1903 & ~n1914;
  assign n1916 = ~n1902 & ~n1915;
  assign n1917 = ~pi058 & pi146;
  assign n1918 = ~pi145 & ~n1917;
  assign n1919 = ~n1916 & n1918;
  assign n1920 = ~pi057 & ~n1919;
  assign n1921 = ~n1916 & ~n1917;
  assign n1922 = pi145 & ~n1921;
  assign n1923 = ~n1920 & ~n1922;
  assign n1924 = ~n1901 & ~n1923;
  assign n1925 = ~n1900 & ~n1924;
  assign n1926 = ~n1899 & ~n1925;
  assign n1927 = ~n1898 & ~n1926;
  assign n1928 = ~n1897 & ~n1927;
  assign n1929 = ~pi055 & pi175;
  assign n1930 = pi055 & ~pi175;
  assign n1931 = ~pi056 & pi176;
  assign n1932 = pi056 & ~pi176;
  assign n1933 = pi058 & ~pi178;
  assign n1934 = ~pi059 & pi179;
  assign n1935 = pi059 & ~pi179;
  assign n1936 = ~pi060 & pi180;
  assign n1937 = pi060 & ~pi180;
  assign n1938 = pi062 & ~pi182;
  assign n1939 = pi061 & ~pi181;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~pi061 & pi181;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = ~n1937 & ~n1942;
  assign n1944 = ~n1936 & ~n1943;
  assign n1945 = ~n1935 & ~n1944;
  assign n1946 = ~n1934 & ~n1945;
  assign n1947 = ~n1933 & ~n1946;
  assign n1948 = ~pi058 & pi178;
  assign n1949 = ~pi177 & ~n1948;
  assign n1950 = ~n1947 & n1949;
  assign n1951 = ~pi057 & ~n1950;
  assign n1952 = ~n1947 & ~n1948;
  assign n1953 = pi177 & ~n1952;
  assign n1954 = ~n1951 & ~n1953;
  assign n1955 = ~n1932 & ~n1954;
  assign n1956 = ~n1931 & ~n1955;
  assign n1957 = ~n1930 & ~n1956;
  assign n1958 = ~n1929 & ~n1957;
  assign n1959 = ~pi055 & pi119;
  assign n1960 = pi055 & ~pi119;
  assign n1961 = ~pi056 & pi120;
  assign n1962 = pi056 & ~pi120;
  assign n1963 = pi058 & ~pi122;
  assign n1964 = ~pi059 & pi123;
  assign n1965 = pi059 & ~pi123;
  assign n1966 = ~pi060 & pi124;
  assign n1967 = pi060 & ~pi124;
  assign n1968 = pi062 & ~pi126;
  assign n1969 = pi061 & ~pi125;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~pi061 & pi125;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1967 & ~n1972;
  assign n1974 = ~n1966 & ~n1973;
  assign n1975 = ~n1965 & ~n1974;
  assign n1976 = ~n1964 & ~n1975;
  assign n1977 = ~n1963 & ~n1976;
  assign n1978 = ~pi058 & pi122;
  assign n1979 = ~pi121 & ~n1978;
  assign n1980 = ~n1977 & n1979;
  assign n1981 = ~pi057 & ~n1980;
  assign n1982 = ~n1977 & ~n1978;
  assign n1983 = pi121 & ~n1982;
  assign n1984 = ~n1981 & ~n1983;
  assign n1985 = ~n1962 & ~n1984;
  assign n1986 = ~n1961 & ~n1985;
  assign n1987 = ~n1960 & ~n1986;
  assign n1988 = ~n1959 & ~n1987;
  assign n1989 = ~n1958 & ~n1988;
  assign n1990 = n1928 & n1989;
  assign n1991 = ~pi055 & pi167;
  assign n1992 = ~pi058 & pi170;
  assign n1993 = pi058 & ~pi170;
  assign n1994 = ~pi059 & pi171;
  assign n1995 = pi059 & ~pi171;
  assign n1996 = ~pi060 & pi172;
  assign n1997 = pi060 & ~pi172;
  assign n1998 = pi062 & ~pi174;
  assign n1999 = pi061 & ~pi173;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~pi061 & pi173;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1997 & ~n2002;
  assign n2004 = ~n1996 & ~n2003;
  assign n2005 = ~n1995 & ~n2004;
  assign n2006 = ~n1994 & ~n2005;
  assign n2007 = ~n1993 & ~n2006;
  assign n2008 = ~n1992 & ~n2007;
  assign n2009 = pi169 & ~n2008;
  assign n2010 = ~pi169 & ~n1992;
  assign n2011 = ~n2007 & n2010;
  assign n2012 = ~pi057 & ~n2011;
  assign n2013 = ~pi056 & pi168;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n2009 & n2014;
  assign n2016 = pi056 & ~pi168;
  assign n2017 = pi055 & ~pi167;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = ~n2015 & n2018;
  assign n2020 = ~n1991 & ~n2019;
  assign n2021 = ~pi055 & pi135;
  assign n2022 = ~pi058 & pi138;
  assign n2023 = pi058 & ~pi138;
  assign n2024 = ~pi059 & pi139;
  assign n2025 = pi059 & ~pi139;
  assign n2026 = ~pi060 & pi140;
  assign n2027 = pi060 & ~pi140;
  assign n2028 = pi062 & ~pi142;
  assign n2029 = pi061 & ~pi141;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = ~pi061 & pi141;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = ~n2027 & ~n2032;
  assign n2034 = ~n2026 & ~n2033;
  assign n2035 = ~n2025 & ~n2034;
  assign n2036 = ~n2024 & ~n2035;
  assign n2037 = ~n2023 & ~n2036;
  assign n2038 = ~n2022 & ~n2037;
  assign n2039 = pi137 & ~n2038;
  assign n2040 = ~pi137 & ~n2022;
  assign n2041 = ~n2037 & n2040;
  assign n2042 = ~pi057 & ~n2041;
  assign n2043 = ~pi056 & pi136;
  assign n2044 = ~n2042 & ~n2043;
  assign n2045 = ~n2039 & n2044;
  assign n2046 = pi056 & ~pi136;
  assign n2047 = pi055 & ~pi135;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~n2045 & n2048;
  assign n2050 = ~n2021 & ~n2049;
  assign n2051 = ~n2020 & ~n2050;
  assign n2052 = ~pi055 & pi127;
  assign n2053 = ~pi058 & pi130;
  assign n2054 = pi058 & ~pi130;
  assign n2055 = ~pi059 & pi131;
  assign n2056 = pi059 & ~pi131;
  assign n2057 = ~pi060 & pi132;
  assign n2058 = pi060 & ~pi132;
  assign n2059 = pi062 & ~pi134;
  assign n2060 = pi061 & ~pi133;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = ~pi061 & pi133;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2058 & ~n2063;
  assign n2065 = ~n2057 & ~n2064;
  assign n2066 = ~n2056 & ~n2065;
  assign n2067 = ~n2055 & ~n2066;
  assign n2068 = ~n2054 & ~n2067;
  assign n2069 = ~n2053 & ~n2068;
  assign n2070 = pi129 & ~n2069;
  assign n2071 = ~pi129 & ~n2053;
  assign n2072 = ~n2068 & n2071;
  assign n2073 = ~pi057 & ~n2072;
  assign n2074 = ~pi056 & pi128;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = ~n2070 & n2075;
  assign n2077 = pi056 & ~pi128;
  assign n2078 = pi055 & ~pi127;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = ~n2076 & n2079;
  assign n2081 = ~n2052 & ~n2080;
  assign n2082 = ~pi055 & pi095;
  assign n2083 = ~pi058 & pi098;
  assign n2084 = pi058 & ~pi098;
  assign n2085 = ~pi059 & pi099;
  assign n2086 = pi059 & ~pi099;
  assign n2087 = ~pi060 & pi100;
  assign n2088 = pi060 & ~pi100;
  assign n2089 = pi062 & ~pi102;
  assign n2090 = pi061 & ~pi101;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~pi061 & pi101;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = ~n2088 & ~n2093;
  assign n2095 = ~n2087 & ~n2094;
  assign n2096 = ~n2086 & ~n2095;
  assign n2097 = ~n2085 & ~n2096;
  assign n2098 = ~n2084 & ~n2097;
  assign n2099 = ~n2083 & ~n2098;
  assign n2100 = ~pi057 & ~n2099;
  assign n2101 = pi057 & ~n2083;
  assign n2102 = ~n2098 & n2101;
  assign n2103 = pi097 & ~n2102;
  assign n2104 = ~pi056 & pi096;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = ~n2100 & n2105;
  assign n2107 = pi056 & ~pi096;
  assign n2108 = pi055 & ~pi095;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~n2106 & n2109;
  assign n2111 = ~n2082 & ~n2110;
  assign n2112 = ~n2081 & ~n2111;
  assign n2113 = n2051 & n2112;
  assign n2114 = ~pi055 & pi207;
  assign n2115 = ~pi058 & pi210;
  assign n2116 = pi058 & ~pi210;
  assign n2117 = ~pi059 & pi211;
  assign n2118 = pi059 & ~pi211;
  assign n2119 = ~pi060 & pi212;
  assign n2120 = pi060 & ~pi212;
  assign n2121 = pi062 & ~pi214;
  assign n2122 = pi061 & ~pi213;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = ~pi061 & pi213;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = ~n2120 & ~n2125;
  assign n2127 = ~n2119 & ~n2126;
  assign n2128 = ~n2118 & ~n2127;
  assign n2129 = ~n2117 & ~n2128;
  assign n2130 = ~n2116 & ~n2129;
  assign n2131 = ~n2115 & ~n2130;
  assign n2132 = pi209 & ~n2131;
  assign n2133 = ~pi209 & ~n2115;
  assign n2134 = ~n2130 & n2133;
  assign n2135 = ~pi057 & ~n2134;
  assign n2136 = ~pi056 & pi208;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2132 & n2137;
  assign n2139 = pi056 & ~pi208;
  assign n2140 = pi055 & ~pi207;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~n2138 & n2141;
  assign n2143 = ~n2114 & ~n2142;
  assign n2144 = pi003 & ~n501;
  assign n2145 = ~n500 & n2144;
  assign n2146 = ~n2143 & n2145;
  assign n2147 = ~pi055 & pi223;
  assign n2148 = ~pi058 & pi226;
  assign n2149 = pi058 & ~pi226;
  assign n2150 = ~pi059 & pi227;
  assign n2151 = pi059 & ~pi227;
  assign n2152 = ~pi060 & pi228;
  assign n2153 = pi060 & ~pi228;
  assign n2154 = pi062 & ~pi230;
  assign n2155 = pi061 & ~pi229;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~pi061 & pi229;
  assign n2158 = ~n2156 & ~n2157;
  assign n2159 = ~n2153 & ~n2158;
  assign n2160 = ~n2152 & ~n2159;
  assign n2161 = ~n2151 & ~n2160;
  assign n2162 = ~n2150 & ~n2161;
  assign n2163 = ~n2149 & ~n2162;
  assign n2164 = ~n2148 & ~n2163;
  assign n2165 = pi225 & ~n2164;
  assign n2166 = ~pi225 & ~n2148;
  assign n2167 = ~n2163 & n2166;
  assign n2168 = ~pi057 & ~n2167;
  assign n2169 = ~pi056 & pi224;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n2165 & n2170;
  assign n2172 = pi056 & ~pi224;
  assign n2173 = pi055 & ~pi223;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n2171 & n2174;
  assign n2176 = ~n2147 & ~n2175;
  assign n2177 = ~pi055 & pi199;
  assign n2178 = ~pi058 & pi202;
  assign n2179 = pi058 & ~pi202;
  assign n2180 = ~pi059 & pi203;
  assign n2181 = pi059 & ~pi203;
  assign n2182 = ~pi060 & pi204;
  assign n2183 = pi060 & ~pi204;
  assign n2184 = pi062 & ~pi206;
  assign n2185 = pi061 & ~pi205;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~pi061 & pi205;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = ~n2183 & ~n2188;
  assign n2190 = ~n2182 & ~n2189;
  assign n2191 = ~n2181 & ~n2190;
  assign n2192 = ~n2180 & ~n2191;
  assign n2193 = ~n2179 & ~n2192;
  assign n2194 = ~n2178 & ~n2193;
  assign n2195 = pi201 & ~n2194;
  assign n2196 = ~pi201 & ~n2178;
  assign n2197 = ~n2193 & n2196;
  assign n2198 = ~pi057 & ~n2197;
  assign n2199 = ~pi056 & pi200;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = ~n2195 & n2200;
  assign n2202 = pi056 & ~pi200;
  assign n2203 = pi055 & ~pi199;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = ~n2201 & n2204;
  assign n2206 = ~n2177 & ~n2205;
  assign n2207 = ~n2176 & ~n2206;
  assign n2208 = n2146 & n2207;
  assign n2209 = n2113 & n2208;
  assign n2210 = n1990 & n2209;
  assign n2211 = n1867 & n2210;
  assign n2212 = n1744 & n2211;
  assign n2213 = ~n1373 & n2212;
  assign n2214 = n564 & ~n595;
  assign n2215 = n844 & n2214;
  assign n2216 = n1362 & n2215;
  assign n2217 = ~n1372 & n2216;
  assign n2218 = pi004 & ~n501;
  assign n2219 = ~n566 & ~n1465;
  assign n2220 = n2218 & n2219;
  assign n2221 = ~n500 & n2220;
  assign n2222 = ~n594 & ~n1493;
  assign n2223 = n2221 & n2222;
  assign n2224 = pi002 & ~n1173;
  assign n2225 = ~n1144 & n2224;
  assign n2226 = ~n1115 & n2225;
  assign n2227 = ~n1086 & n2226;
  assign n2228 = n1057 & n2227;
  assign n2229 = n1239 & n2228;
  assign n2230 = n1360 & n2229;
  assign n2231 = n968 & n2230;
  assign n2232 = n845 & n2231;
  assign n2233 = ~n2223 & ~n2232;
  assign n2234 = ~n2217 & n2233;
  assign po002 = n2213 | ~n2234;
  assign n2236 = po144 & ~n2143;
  assign n2237 = n2207 & n2236;
  assign n2238 = n2113 & n2237;
  assign n2239 = n1990 & n2238;
  assign n2240 = n1867 & n2239;
  assign n2241 = n1744 & n2240;
  assign n2242 = ~n1373 & n2241;
  assign n2243 = n1371 & n2215;
  assign n2244 = n1373 & ~n2243;
  assign n2245 = ~po144 & ~n1372;
  assign n2246 = ~n501 & ~n566;
  assign n2247 = ~n1465 & n2246;
  assign n2248 = ~n500 & n2247;
  assign po145 = n2222 & n2248;
  assign n2250 = n1494 & ~po145;
  assign n2251 = n1434 & ~n1464;
  assign n2252 = ~n2250 & n2251;
  assign n2253 = n1743 & n2252;
  assign n2254 = pi003 & ~n2143;
  assign n2255 = n2207 & n2254;
  assign n2256 = n2113 & n2255;
  assign n2257 = n1990 & n2256;
  assign n2258 = n1867 & n2257;
  assign n2259 = n2253 & n2258;
  assign n2260 = ~n2245 & n2259;
  assign n2261 = ~n2244 & n2260;
  assign n2262 = ~n2242 & n2261;
  assign n2263 = n936 & ~n2241;
  assign n2264 = n595 & ~po145;
  assign n2265 = n564 & n719;
  assign n2266 = n658 & n842;
  assign n2267 = n2265 & n2266;
  assign n2268 = ~n2264 & n2267;
  assign n2269 = ~n875 & ~n1270;
  assign n2270 = ~n905 & ~n966;
  assign n2271 = n2269 & n2270;
  assign n2272 = n781 & n1239;
  assign n2273 = n1178 & n1359;
  assign n2274 = n2272 & n2273;
  assign n2275 = n2271 & n2274;
  assign n2276 = n2268 & n2275;
  assign n2277 = ~n1372 & n2276;
  assign n2278 = ~n2243 & n2277;
  assign n2279 = ~n2263 & n2278;
  assign n2280 = pi073 & ~pi081;
  assign n2281 = ~pi074 & pi082;
  assign n2282 = pi074 & ~pi082;
  assign n2283 = ~pi075 & pi083;
  assign n2284 = pi075 & ~pi083;
  assign n2285 = ~pi076 & pi084;
  assign n2286 = pi076 & ~pi084;
  assign n2287 = pi078 & ~pi086;
  assign n2288 = pi077 & ~pi085;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = ~pi077 & pi085;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n2286 & ~n2291;
  assign n2293 = ~n2285 & ~n2292;
  assign n2294 = ~n2284 & ~n2293;
  assign n2295 = ~n2283 & ~n2294;
  assign n2296 = ~n2282 & ~n2295;
  assign n2297 = ~n2281 & ~n2296;
  assign n2298 = ~n2280 & ~n2297;
  assign n2299 = ~pi073 & pi081;
  assign n2300 = ~pi072 & pi080;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = pi071 & ~pi079;
  assign n2304 = pi072 & ~pi080;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n2302 & n2305;
  assign n2307 = ~pi071 & pi079;
  assign n2308 = ~n1435 & ~n1465;
  assign n2309 = ~n2307 & n2308;
  assign n2310 = pi006 & ~n501;
  assign n2311 = ~n504 & ~n566;
  assign n2312 = n2310 & n2311;
  assign n2313 = n2309 & n2312;
  assign n2314 = ~n2306 & n2313;
  assign n2315 = ~n500 & n2314;
  assign n2316 = ~n532 & ~n594;
  assign n2317 = ~n1463 & ~n1493;
  assign n2318 = n2316 & n2317;
  assign n2319 = n2315 & n2318;
  assign n2320 = ~n2279 & ~n2319;
  assign n2321 = ~n2262 & n2320;
  assign n2322 = ~n1494 & ~n2242;
  assign n2323 = ~n595 & ~n1372;
  assign n2324 = ~n2243 & n2323;
  assign n2325 = pi004 & ~po145;
  assign n2326 = ~n2245 & n2325;
  assign n2327 = ~n2324 & n2326;
  assign n2328 = ~n2322 & n2327;
  assign n2329 = ~n1774 & ~n2242;
  assign n2330 = ~n905 & ~n1372;
  assign n2331 = ~n2243 & n2330;
  assign n2332 = pi005 & ~n501;
  assign n2333 = n2219 & n2332;
  assign n2334 = ~n500 & n2333;
  assign n2335 = ~pi071 & pi135;
  assign n2336 = pi073 & ~pi137;
  assign n2337 = ~pi074 & pi138;
  assign n2338 = pi074 & ~pi138;
  assign n2339 = ~pi075 & pi139;
  assign n2340 = pi075 & ~pi139;
  assign n2341 = ~pi076 & pi140;
  assign n2342 = pi076 & ~pi140;
  assign n2343 = pi078 & ~pi142;
  assign n2344 = pi077 & ~pi141;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~pi077 & pi141;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n2342 & ~n2347;
  assign n2349 = ~n2341 & ~n2348;
  assign n2350 = ~n2340 & ~n2349;
  assign n2351 = ~n2339 & ~n2350;
  assign n2352 = ~n2338 & ~n2351;
  assign n2353 = ~n2337 & ~n2352;
  assign n2354 = ~n2336 & ~n2353;
  assign n2355 = ~pi073 & pi137;
  assign n2356 = ~pi072 & pi136;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = ~n2354 & n2357;
  assign n2359 = pi071 & ~pi135;
  assign n2360 = pi072 & ~pi136;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n2358 & n2361;
  assign n2363 = ~n2335 & ~n2362;
  assign n2364 = ~pi071 & pi095;
  assign n2365 = pi073 & ~pi097;
  assign n2366 = ~pi074 & pi098;
  assign n2367 = pi074 & ~pi098;
  assign n2368 = ~pi075 & pi099;
  assign n2369 = pi075 & ~pi099;
  assign n2370 = ~pi076 & pi100;
  assign n2371 = pi076 & ~pi100;
  assign n2372 = pi078 & ~pi102;
  assign n2373 = pi077 & ~pi101;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~pi077 & pi101;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n2371 & ~n2376;
  assign n2378 = ~n2370 & ~n2377;
  assign n2379 = ~n2369 & ~n2378;
  assign n2380 = ~n2368 & ~n2379;
  assign n2381 = ~n2367 & ~n2380;
  assign n2382 = ~n2366 & ~n2381;
  assign n2383 = ~n2365 & ~n2382;
  assign n2384 = ~pi073 & pi097;
  assign n2385 = ~pi072 & pi096;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2383 & n2386;
  assign n2388 = pi071 & ~pi095;
  assign n2389 = pi072 & ~pi096;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n2387 & n2390;
  assign n2392 = ~n2364 & ~n2391;
  assign n2393 = ~n2363 & ~n2392;
  assign n2394 = n2222 & n2393;
  assign n2395 = n2334 & n2394;
  assign n2396 = ~pi071 & pi239;
  assign n2397 = pi073 & ~pi241;
  assign n2398 = ~pi074 & pi242;
  assign n2399 = pi074 & ~pi242;
  assign n2400 = ~pi075 & pi243;
  assign n2401 = pi075 & ~pi243;
  assign n2402 = ~pi076 & pi244;
  assign n2403 = pi076 & ~pi244;
  assign n2404 = pi078 & ~pi246;
  assign n2405 = pi077 & ~pi245;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~pi077 & pi245;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = ~n2403 & ~n2408;
  assign n2410 = ~n2402 & ~n2409;
  assign n2411 = ~n2401 & ~n2410;
  assign n2412 = ~n2400 & ~n2411;
  assign n2413 = ~n2399 & ~n2412;
  assign n2414 = ~n2398 & ~n2413;
  assign n2415 = ~n2397 & ~n2414;
  assign n2416 = ~pi073 & pi241;
  assign n2417 = ~pi072 & pi240;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = ~n2415 & n2418;
  assign n2420 = pi071 & ~pi239;
  assign n2421 = pi072 & ~pi240;
  assign n2422 = ~n2420 & ~n2421;
  assign n2423 = ~n2419 & n2422;
  assign n2424 = ~n2396 & ~n2423;
  assign n2425 = ~pi071 & pi183;
  assign n2426 = pi073 & ~pi185;
  assign n2427 = ~pi074 & pi186;
  assign n2428 = pi074 & ~pi186;
  assign n2429 = ~pi075 & pi187;
  assign n2430 = pi075 & ~pi187;
  assign n2431 = ~pi076 & pi188;
  assign n2432 = pi076 & ~pi188;
  assign n2433 = pi078 & ~pi190;
  assign n2434 = pi077 & ~pi189;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = ~pi077 & pi189;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2432 & ~n2437;
  assign n2439 = ~n2431 & ~n2438;
  assign n2440 = ~n2430 & ~n2439;
  assign n2441 = ~n2429 & ~n2440;
  assign n2442 = ~n2428 & ~n2441;
  assign n2443 = ~n2427 & ~n2442;
  assign n2444 = ~n2426 & ~n2443;
  assign n2445 = ~pi073 & pi185;
  assign n2446 = ~pi072 & pi184;
  assign n2447 = ~n2445 & ~n2446;
  assign n2448 = ~n2444 & n2447;
  assign n2449 = pi071 & ~pi183;
  assign n2450 = pi072 & ~pi184;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = ~n2448 & n2451;
  assign n2453 = ~n2425 & ~n2452;
  assign n2454 = ~n2424 & ~n2453;
  assign n2455 = ~pi071 & pi199;
  assign n2456 = pi073 & ~pi201;
  assign n2457 = ~pi074 & pi202;
  assign n2458 = pi074 & ~pi202;
  assign n2459 = ~pi075 & pi203;
  assign n2460 = pi075 & ~pi203;
  assign n2461 = ~pi076 & pi204;
  assign n2462 = pi076 & ~pi204;
  assign n2463 = pi078 & ~pi206;
  assign n2464 = pi077 & ~pi205;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~pi077 & pi205;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n2462 & ~n2467;
  assign n2469 = ~n2461 & ~n2468;
  assign n2470 = ~n2460 & ~n2469;
  assign n2471 = ~n2459 & ~n2470;
  assign n2472 = ~n2458 & ~n2471;
  assign n2473 = ~n2457 & ~n2472;
  assign n2474 = ~n2456 & ~n2473;
  assign n2475 = ~pi073 & pi201;
  assign n2476 = ~pi072 & pi200;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2474 & n2477;
  assign n2479 = pi071 & ~pi199;
  assign n2480 = pi072 & ~pi200;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = ~n2478 & n2481;
  assign n2483 = ~n2455 & ~n2482;
  assign n2484 = ~pi071 & pi207;
  assign n2485 = pi073 & ~pi209;
  assign n2486 = ~pi074 & pi210;
  assign n2487 = pi074 & ~pi210;
  assign n2488 = ~pi075 & pi211;
  assign n2489 = pi075 & ~pi211;
  assign n2490 = ~pi076 & pi212;
  assign n2491 = pi076 & ~pi212;
  assign n2492 = pi078 & ~pi214;
  assign n2493 = pi077 & ~pi213;
  assign n2494 = ~n2492 & ~n2493;
  assign n2495 = ~pi077 & pi213;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = ~n2491 & ~n2496;
  assign n2498 = ~n2490 & ~n2497;
  assign n2499 = ~n2489 & ~n2498;
  assign n2500 = ~n2488 & ~n2499;
  assign n2501 = ~n2487 & ~n2500;
  assign n2502 = ~n2486 & ~n2501;
  assign n2503 = ~n2485 & ~n2502;
  assign n2504 = ~pi073 & pi209;
  assign n2505 = ~pi072 & pi208;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = ~n2503 & n2506;
  assign n2508 = pi071 & ~pi207;
  assign n2509 = pi072 & ~pi208;
  assign n2510 = ~n2508 & ~n2509;
  assign n2511 = ~n2507 & n2510;
  assign n2512 = ~n2484 & ~n2511;
  assign n2513 = ~n2483 & ~n2512;
  assign n2514 = n2454 & n2513;
  assign n2515 = ~pi071 & pi255;
  assign n2516 = pi073 & ~pi257;
  assign n2517 = ~pi074 & pi258;
  assign n2518 = pi074 & ~pi258;
  assign n2519 = ~pi075 & pi259;
  assign n2520 = pi075 & ~pi259;
  assign n2521 = ~pi076 & pi260;
  assign n2522 = pi076 & ~pi260;
  assign n2523 = pi078 & ~pi262;
  assign n2524 = pi077 & ~pi261;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = ~pi077 & pi261;
  assign n2527 = ~n2525 & ~n2526;
  assign n2528 = ~n2522 & ~n2527;
  assign n2529 = ~n2521 & ~n2528;
  assign n2530 = ~n2520 & ~n2529;
  assign n2531 = ~n2519 & ~n2530;
  assign n2532 = ~n2518 & ~n2531;
  assign n2533 = ~n2517 & ~n2532;
  assign n2534 = ~n2516 & ~n2533;
  assign n2535 = ~pi073 & pi257;
  assign n2536 = ~pi072 & pi256;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = ~n2534 & n2537;
  assign n2539 = pi071 & ~pi255;
  assign n2540 = pi072 & ~pi256;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~n2538 & n2541;
  assign n2543 = ~n2515 & ~n2542;
  assign n2544 = ~pi071 & pi247;
  assign n2545 = pi073 & ~pi249;
  assign n2546 = ~pi074 & pi250;
  assign n2547 = pi074 & ~pi250;
  assign n2548 = ~pi075 & pi251;
  assign n2549 = pi075 & ~pi251;
  assign n2550 = ~pi076 & pi252;
  assign n2551 = pi076 & ~pi252;
  assign n2552 = pi078 & ~pi254;
  assign n2553 = pi077 & ~pi253;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~pi077 & pi253;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2551 & ~n2556;
  assign n2558 = ~n2550 & ~n2557;
  assign n2559 = ~n2549 & ~n2558;
  assign n2560 = ~n2548 & ~n2559;
  assign n2561 = ~n2547 & ~n2560;
  assign n2562 = ~n2546 & ~n2561;
  assign n2563 = ~n2545 & ~n2562;
  assign n2564 = ~pi073 & pi249;
  assign n2565 = ~pi072 & pi248;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = ~n2563 & n2566;
  assign n2568 = pi071 & ~pi247;
  assign n2569 = pi072 & ~pi248;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2567 & n2570;
  assign n2572 = ~n2544 & ~n2571;
  assign n2573 = ~n2543 & ~n2572;
  assign n2574 = ~pi071 & pi263;
  assign n2575 = pi073 & ~pi265;
  assign n2576 = ~pi074 & pi266;
  assign n2577 = pi074 & ~pi266;
  assign n2578 = ~pi075 & pi267;
  assign n2579 = pi075 & ~pi267;
  assign n2580 = ~pi076 & pi268;
  assign n2581 = pi076 & ~pi268;
  assign n2582 = pi078 & ~pi270;
  assign n2583 = pi077 & ~pi269;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = ~pi077 & pi269;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2581 & ~n2586;
  assign n2588 = ~n2580 & ~n2587;
  assign n2589 = ~n2579 & ~n2588;
  assign n2590 = ~n2578 & ~n2589;
  assign n2591 = ~n2577 & ~n2590;
  assign n2592 = ~n2576 & ~n2591;
  assign n2593 = ~n2575 & ~n2592;
  assign n2594 = ~pi073 & pi265;
  assign n2595 = ~pi072 & pi264;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = ~n2593 & n2596;
  assign n2598 = pi071 & ~pi263;
  assign n2599 = pi072 & ~pi264;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = ~n2597 & n2600;
  assign n2602 = ~n2574 & ~n2601;
  assign n2603 = ~pi071 & pi231;
  assign n2604 = pi073 & ~pi233;
  assign n2605 = ~pi074 & pi234;
  assign n2606 = pi074 & ~pi234;
  assign n2607 = ~pi075 & pi235;
  assign n2608 = pi075 & ~pi235;
  assign n2609 = ~pi076 & pi236;
  assign n2610 = pi076 & ~pi236;
  assign n2611 = pi078 & ~pi238;
  assign n2612 = pi077 & ~pi237;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~pi077 & pi237;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = ~n2610 & ~n2615;
  assign n2617 = ~n2609 & ~n2616;
  assign n2618 = ~n2608 & ~n2617;
  assign n2619 = ~n2607 & ~n2618;
  assign n2620 = ~n2606 & ~n2619;
  assign n2621 = ~n2605 & ~n2620;
  assign n2622 = ~n2604 & ~n2621;
  assign n2623 = ~pi073 & pi233;
  assign n2624 = ~pi072 & pi232;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = ~n2622 & n2625;
  assign n2627 = pi071 & ~pi231;
  assign n2628 = pi072 & ~pi232;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2626 & n2629;
  assign n2631 = ~n2603 & ~n2630;
  assign n2632 = ~n2602 & ~n2631;
  assign n2633 = n2573 & n2632;
  assign n2634 = n2514 & n2633;
  assign n2635 = ~pi071 & pi223;
  assign n2636 = pi073 & ~pi225;
  assign n2637 = ~pi074 & pi226;
  assign n2638 = pi074 & ~pi226;
  assign n2639 = ~pi075 & pi227;
  assign n2640 = pi075 & ~pi227;
  assign n2641 = ~pi076 & pi228;
  assign n2642 = pi076 & ~pi228;
  assign n2643 = pi078 & ~pi230;
  assign n2644 = pi077 & ~pi229;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = ~pi077 & pi229;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = ~n2642 & ~n2647;
  assign n2649 = ~n2641 & ~n2648;
  assign n2650 = ~n2640 & ~n2649;
  assign n2651 = ~n2639 & ~n2650;
  assign n2652 = ~n2638 & ~n2651;
  assign n2653 = ~n2637 & ~n2652;
  assign n2654 = ~n2636 & ~n2653;
  assign n2655 = ~pi073 & pi225;
  assign n2656 = ~pi072 & pi224;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = ~n2654 & n2657;
  assign n2659 = pi071 & ~pi223;
  assign n2660 = pi072 & ~pi224;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2658 & n2661;
  assign n2663 = ~n2635 & ~n2662;
  assign n2664 = ~pi071 & pi111;
  assign n2665 = pi073 & ~pi113;
  assign n2666 = ~pi074 & pi114;
  assign n2667 = pi074 & ~pi114;
  assign n2668 = ~pi075 & pi115;
  assign n2669 = pi075 & ~pi115;
  assign n2670 = ~pi076 & pi116;
  assign n2671 = pi076 & ~pi116;
  assign n2672 = pi078 & ~pi118;
  assign n2673 = pi077 & ~pi117;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = ~pi077 & pi117;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2671 & ~n2676;
  assign n2678 = ~n2670 & ~n2677;
  assign n2679 = ~n2669 & ~n2678;
  assign n2680 = ~n2668 & ~n2679;
  assign n2681 = ~n2667 & ~n2680;
  assign n2682 = ~n2666 & ~n2681;
  assign n2683 = ~n2665 & ~n2682;
  assign n2684 = ~pi073 & pi113;
  assign n2685 = ~pi072 & pi112;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = ~n2683 & n2686;
  assign n2688 = pi071 & ~pi111;
  assign n2689 = pi072 & ~pi112;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = ~n2687 & n2690;
  assign n2692 = ~n2664 & ~n2691;
  assign n2693 = ~n2663 & ~n2692;
  assign n2694 = ~pi071 & pi127;
  assign n2695 = pi073 & ~pi129;
  assign n2696 = ~pi074 & pi130;
  assign n2697 = pi074 & ~pi130;
  assign n2698 = ~pi075 & pi131;
  assign n2699 = pi075 & ~pi131;
  assign n2700 = ~pi076 & pi132;
  assign n2701 = pi076 & ~pi132;
  assign n2702 = pi078 & ~pi134;
  assign n2703 = pi077 & ~pi133;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~pi077 & pi133;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2701 & ~n2706;
  assign n2708 = ~n2700 & ~n2707;
  assign n2709 = ~n2699 & ~n2708;
  assign n2710 = ~n2698 & ~n2709;
  assign n2711 = ~n2697 & ~n2710;
  assign n2712 = ~n2696 & ~n2711;
  assign n2713 = ~n2695 & ~n2712;
  assign n2714 = ~pi073 & pi129;
  assign n2715 = ~pi072 & pi128;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2713 & n2716;
  assign n2718 = pi071 & ~pi127;
  assign n2719 = pi072 & ~pi128;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = ~n2717 & n2720;
  assign n2722 = ~n2694 & ~n2721;
  assign n2723 = ~n2306 & ~n2307;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2693 & n2724;
  assign n2726 = ~pi071 & pi215;
  assign n2727 = pi073 & ~pi217;
  assign n2728 = ~pi074 & pi218;
  assign n2729 = pi074 & ~pi218;
  assign n2730 = ~pi075 & pi219;
  assign n2731 = pi075 & ~pi219;
  assign n2732 = ~pi076 & pi220;
  assign n2733 = pi076 & ~pi220;
  assign n2734 = pi078 & ~pi222;
  assign n2735 = pi077 & ~pi221;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = ~pi077 & pi221;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = ~n2733 & ~n2738;
  assign n2740 = ~n2732 & ~n2739;
  assign n2741 = ~n2731 & ~n2740;
  assign n2742 = ~n2730 & ~n2741;
  assign n2743 = ~n2729 & ~n2742;
  assign n2744 = ~n2728 & ~n2743;
  assign n2745 = ~n2727 & ~n2744;
  assign n2746 = ~pi073 & pi217;
  assign n2747 = ~pi072 & pi216;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = ~n2745 & n2748;
  assign n2750 = pi071 & ~pi215;
  assign n2751 = pi072 & ~pi216;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = ~n2749 & n2752;
  assign n2754 = ~n2726 & ~n2753;
  assign n2755 = ~pi071 & pi271;
  assign n2756 = pi073 & ~pi273;
  assign n2757 = ~pi074 & pi274;
  assign n2758 = pi074 & ~pi274;
  assign n2759 = ~pi075 & pi275;
  assign n2760 = pi075 & ~pi275;
  assign n2761 = ~pi076 & pi276;
  assign n2762 = pi076 & ~pi276;
  assign n2763 = pi078 & ~pi278;
  assign n2764 = pi077 & ~pi277;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = ~pi077 & pi277;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = ~n2762 & ~n2767;
  assign n2769 = ~n2761 & ~n2768;
  assign n2770 = ~n2760 & ~n2769;
  assign n2771 = ~n2759 & ~n2770;
  assign n2772 = ~n2758 & ~n2771;
  assign n2773 = ~n2757 & ~n2772;
  assign n2774 = ~n2756 & ~n2773;
  assign n2775 = ~pi073 & pi273;
  assign n2776 = ~pi072 & pi272;
  assign n2777 = ~n2775 & ~n2776;
  assign n2778 = ~n2774 & n2777;
  assign n2779 = pi071 & ~pi271;
  assign n2780 = pi072 & ~pi272;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2778 & n2781;
  assign n2783 = ~n2755 & ~n2782;
  assign n2784 = ~n2754 & ~n2783;
  assign n2785 = ~pi071 & pi151;
  assign n2786 = pi073 & ~pi153;
  assign n2787 = ~pi074 & pi154;
  assign n2788 = pi074 & ~pi154;
  assign n2789 = ~pi075 & pi155;
  assign n2790 = pi075 & ~pi155;
  assign n2791 = ~pi076 & pi156;
  assign n2792 = pi076 & ~pi156;
  assign n2793 = pi078 & ~pi158;
  assign n2794 = pi077 & ~pi157;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~pi077 & pi157;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = ~n2792 & ~n2797;
  assign n2799 = ~n2791 & ~n2798;
  assign n2800 = ~n2790 & ~n2799;
  assign n2801 = ~n2789 & ~n2800;
  assign n2802 = ~n2788 & ~n2801;
  assign n2803 = ~n2787 & ~n2802;
  assign n2804 = ~n2786 & ~n2803;
  assign n2805 = ~pi073 & pi153;
  assign n2806 = ~pi072 & pi152;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = ~n2804 & n2807;
  assign n2809 = pi071 & ~pi151;
  assign n2810 = pi072 & ~pi152;
  assign n2811 = ~n2809 & ~n2810;
  assign n2812 = ~n2808 & n2811;
  assign n2813 = ~n2785 & ~n2812;
  assign n2814 = ~pi071 & pi167;
  assign n2815 = pi073 & ~pi169;
  assign n2816 = ~pi074 & pi170;
  assign n2817 = pi074 & ~pi170;
  assign n2818 = ~pi075 & pi171;
  assign n2819 = pi075 & ~pi171;
  assign n2820 = ~pi076 & pi172;
  assign n2821 = pi076 & ~pi172;
  assign n2822 = pi078 & ~pi174;
  assign n2823 = pi077 & ~pi173;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~pi077 & pi173;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = ~n2821 & ~n2826;
  assign n2828 = ~n2820 & ~n2827;
  assign n2829 = ~n2819 & ~n2828;
  assign n2830 = ~n2818 & ~n2829;
  assign n2831 = ~n2817 & ~n2830;
  assign n2832 = ~n2816 & ~n2831;
  assign n2833 = ~n2815 & ~n2832;
  assign n2834 = ~pi073 & pi169;
  assign n2835 = ~pi072 & pi168;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = ~n2833 & n2836;
  assign n2838 = pi071 & ~pi167;
  assign n2839 = pi072 & ~pi168;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = ~n2837 & n2840;
  assign n2842 = ~n2814 & ~n2841;
  assign n2843 = ~n2813 & ~n2842;
  assign n2844 = n2784 & n2843;
  assign n2845 = n2725 & n2844;
  assign n2846 = n2634 & n2845;
  assign n2847 = n2395 & n2846;
  assign n2848 = ~pi071 & pi119;
  assign n2849 = pi071 & ~pi119;
  assign n2850 = ~pi072 & pi120;
  assign n2851 = pi072 & ~pi120;
  assign n2852 = ~pi073 & pi121;
  assign n2853 = pi073 & ~pi121;
  assign n2854 = ~pi074 & pi122;
  assign n2855 = pi074 & ~pi122;
  assign n2856 = ~pi075 & pi123;
  assign n2857 = pi075 & ~pi123;
  assign n2858 = ~pi076 & pi124;
  assign n2859 = pi076 & ~pi124;
  assign n2860 = pi078 & ~pi126;
  assign n2861 = pi077 & ~pi125;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = ~pi077 & pi125;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = ~n2859 & ~n2864;
  assign n2866 = ~n2858 & ~n2865;
  assign n2867 = ~n2857 & ~n2866;
  assign n2868 = ~n2856 & ~n2867;
  assign n2869 = ~n2855 & ~n2868;
  assign n2870 = ~n2854 & ~n2869;
  assign n2871 = ~n2853 & ~n2870;
  assign n2872 = ~n2852 & ~n2871;
  assign n2873 = ~n2851 & ~n2872;
  assign n2874 = ~n2850 & ~n2873;
  assign n2875 = ~n2849 & ~n2874;
  assign n2876 = ~n2848 & ~n2875;
  assign n2877 = ~pi071 & pi103;
  assign n2878 = pi071 & ~pi103;
  assign n2879 = ~pi072 & pi104;
  assign n2880 = pi072 & ~pi104;
  assign n2881 = ~pi073 & pi105;
  assign n2882 = pi073 & ~pi105;
  assign n2883 = ~pi074 & pi106;
  assign n2884 = pi074 & ~pi106;
  assign n2885 = ~pi075 & pi107;
  assign n2886 = pi075 & ~pi107;
  assign n2887 = ~pi076 & pi108;
  assign n2888 = pi076 & ~pi108;
  assign n2889 = pi078 & ~pi110;
  assign n2890 = pi077 & ~pi109;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = ~pi077 & pi109;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = ~n2888 & ~n2893;
  assign n2895 = ~n2887 & ~n2894;
  assign n2896 = ~n2886 & ~n2895;
  assign n2897 = ~n2885 & ~n2896;
  assign n2898 = ~n2884 & ~n2897;
  assign n2899 = ~n2883 & ~n2898;
  assign n2900 = ~n2882 & ~n2899;
  assign n2901 = ~n2881 & ~n2900;
  assign n2902 = ~n2880 & ~n2901;
  assign n2903 = ~n2879 & ~n2902;
  assign n2904 = ~n2878 & ~n2903;
  assign n2905 = ~n2877 & ~n2904;
  assign n2906 = ~pi071 & pi175;
  assign n2907 = pi071 & ~pi175;
  assign n2908 = ~pi072 & pi176;
  assign n2909 = pi072 & ~pi176;
  assign n2910 = ~pi073 & pi177;
  assign n2911 = pi073 & ~pi177;
  assign n2912 = ~pi074 & pi178;
  assign n2913 = pi074 & ~pi178;
  assign n2914 = ~pi075 & pi179;
  assign n2915 = pi075 & ~pi179;
  assign n2916 = ~pi076 & pi180;
  assign n2917 = pi076 & ~pi180;
  assign n2918 = pi078 & ~pi182;
  assign n2919 = pi077 & ~pi181;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = ~pi077 & pi181;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = ~n2917 & ~n2922;
  assign n2924 = ~n2916 & ~n2923;
  assign n2925 = ~n2915 & ~n2924;
  assign n2926 = ~n2914 & ~n2925;
  assign n2927 = ~n2913 & ~n2926;
  assign n2928 = ~n2912 & ~n2927;
  assign n2929 = ~n2911 & ~n2928;
  assign n2930 = ~n2910 & ~n2929;
  assign n2931 = ~n2909 & ~n2930;
  assign n2932 = ~n2908 & ~n2931;
  assign n2933 = ~n2907 & ~n2932;
  assign n2934 = ~n2906 & ~n2933;
  assign n2935 = ~n2905 & ~n2934;
  assign n2936 = ~n2876 & n2935;
  assign n2937 = ~pi071 & pi143;
  assign n2938 = pi071 & ~pi143;
  assign n2939 = ~pi072 & pi144;
  assign n2940 = pi072 & ~pi144;
  assign n2941 = ~pi073 & pi145;
  assign n2942 = pi073 & ~pi145;
  assign n2943 = ~pi074 & pi146;
  assign n2944 = pi074 & ~pi146;
  assign n2945 = ~pi075 & pi147;
  assign n2946 = pi075 & ~pi147;
  assign n2947 = ~pi076 & pi148;
  assign n2948 = pi076 & ~pi148;
  assign n2949 = pi078 & ~pi150;
  assign n2950 = pi077 & ~pi149;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~pi077 & pi149;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~n2948 & ~n2953;
  assign n2955 = ~n2947 & ~n2954;
  assign n2956 = ~n2946 & ~n2955;
  assign n2957 = ~n2945 & ~n2956;
  assign n2958 = ~n2944 & ~n2957;
  assign n2959 = ~n2943 & ~n2958;
  assign n2960 = ~n2942 & ~n2959;
  assign n2961 = ~n2941 & ~n2960;
  assign n2962 = ~n2940 & ~n2961;
  assign n2963 = ~n2939 & ~n2962;
  assign n2964 = ~n2938 & ~n2963;
  assign n2965 = ~n2937 & ~n2964;
  assign n2966 = ~pi071 & pi087;
  assign n2967 = pi071 & ~pi087;
  assign n2968 = ~pi072 & pi088;
  assign n2969 = pi072 & ~pi088;
  assign n2970 = ~pi073 & pi089;
  assign n2971 = pi073 & ~pi089;
  assign n2972 = ~pi074 & pi090;
  assign n2973 = pi074 & ~pi090;
  assign n2974 = ~pi075 & pi091;
  assign n2975 = pi075 & ~pi091;
  assign n2976 = ~pi076 & pi092;
  assign n2977 = pi076 & ~pi092;
  assign n2978 = pi078 & ~pi094;
  assign n2979 = pi077 & ~pi093;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~pi077 & pi093;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2977 & ~n2982;
  assign n2984 = ~n2976 & ~n2983;
  assign n2985 = ~n2975 & ~n2984;
  assign n2986 = ~n2974 & ~n2985;
  assign n2987 = ~n2973 & ~n2986;
  assign n2988 = ~n2972 & ~n2987;
  assign n2989 = ~n2971 & ~n2988;
  assign n2990 = ~n2970 & ~n2989;
  assign n2991 = ~n2969 & ~n2990;
  assign n2992 = ~n2968 & ~n2991;
  assign n2993 = ~n2967 & ~n2992;
  assign n2994 = ~n2966 & ~n2993;
  assign n2995 = ~n2965 & ~n2994;
  assign n2996 = ~pi071 & pi191;
  assign n2997 = pi071 & ~pi191;
  assign n2998 = ~pi072 & pi192;
  assign n2999 = pi072 & ~pi192;
  assign n3000 = ~pi073 & pi193;
  assign n3001 = pi073 & ~pi193;
  assign n3002 = ~pi074 & pi194;
  assign n3003 = pi074 & ~pi194;
  assign n3004 = ~pi075 & pi195;
  assign n3005 = pi075 & ~pi195;
  assign n3006 = ~pi076 & pi196;
  assign n3007 = pi076 & ~pi196;
  assign n3008 = pi078 & ~pi198;
  assign n3009 = pi077 & ~pi197;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = ~pi077 & pi197;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n3007 & ~n3012;
  assign n3014 = ~n3006 & ~n3013;
  assign n3015 = ~n3005 & ~n3014;
  assign n3016 = ~n3004 & ~n3015;
  assign n3017 = ~n3003 & ~n3016;
  assign n3018 = ~n3002 & ~n3017;
  assign n3019 = ~n3001 & ~n3018;
  assign n3020 = ~n3000 & ~n3019;
  assign n3021 = ~n2999 & ~n3020;
  assign n3022 = ~n2998 & ~n3021;
  assign n3023 = ~n2997 & ~n3022;
  assign n3024 = ~n2996 & ~n3023;
  assign n3025 = ~pi071 & pi159;
  assign n3026 = pi071 & ~pi159;
  assign n3027 = ~pi072 & pi160;
  assign n3028 = pi072 & ~pi160;
  assign n3029 = ~pi073 & pi161;
  assign n3030 = pi073 & ~pi161;
  assign n3031 = ~pi074 & pi162;
  assign n3032 = pi074 & ~pi162;
  assign n3033 = ~pi075 & pi163;
  assign n3034 = pi075 & ~pi163;
  assign n3035 = ~pi076 & pi164;
  assign n3036 = pi076 & ~pi164;
  assign n3037 = pi078 & ~pi166;
  assign n3038 = pi077 & ~pi165;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = ~pi077 & pi165;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3036 & ~n3041;
  assign n3043 = ~n3035 & ~n3042;
  assign n3044 = ~n3034 & ~n3043;
  assign n3045 = ~n3033 & ~n3044;
  assign n3046 = ~n3032 & ~n3045;
  assign n3047 = ~n3031 & ~n3046;
  assign n3048 = ~n3030 & ~n3047;
  assign n3049 = ~n3029 & ~n3048;
  assign n3050 = ~n3028 & ~n3049;
  assign n3051 = ~n3027 & ~n3050;
  assign n3052 = ~n3026 & ~n3051;
  assign n3053 = ~n3025 & ~n3052;
  assign n3054 = ~n3024 & ~n3053;
  assign n3055 = n2995 & n3054;
  assign n3056 = n2936 & n3055;
  assign n3057 = n2847 & n3056;
  assign n3058 = ~n2331 & n3057;
  assign n3059 = ~n2329 & n3058;
  assign n3060 = ~n2328 & ~n3059;
  assign po003 = ~n2321 | ~n3060;
  assign n3062 = n2248 & n2394;
  assign n3063 = n2846 & n3062;
  assign n3064 = n3056 & n3063;
  assign n3065 = ~n2331 & n3064;
  assign n3066 = ~n2329 & n3065;
  assign n3067 = ~n2994 & ~n3066;
  assign n3068 = ~n1526 & ~n1740;
  assign n3069 = ~n1556 & ~n1587;
  assign n3070 = n3068 & n3069;
  assign n3071 = ~n1649 & ~n2111;
  assign n3072 = ~n1679 & ~n1710;
  assign n3073 = n3071 & n3072;
  assign n3074 = n3070 & n3073;
  assign n3075 = ~n1403 & ~n1617;
  assign n3076 = ~n1433 & ~n1464;
  assign n3077 = n3075 & n3076;
  assign n3078 = ~n2250 & n3077;
  assign n3079 = n3074 & n3078;
  assign n3080 = ~n1804 & ~n1835;
  assign n3081 = ~n1865 & n3080;
  assign n3082 = ~n1927 & ~n1958;
  assign n3083 = ~n1774 & ~n1988;
  assign n3084 = n3082 & n3083;
  assign n3085 = ~n2020 & ~n2206;
  assign n3086 = ~n2050 & ~n2081;
  assign n3087 = n3085 & n3086;
  assign n3088 = ~n2143 & ~n2176;
  assign n3089 = ~n1897 & n3088;
  assign n3090 = n3087 & n3089;
  assign n3091 = n3084 & n3090;
  assign n3092 = n3081 & n3091;
  assign n3093 = n3079 & n3092;
  assign n3094 = ~n2245 & n3093;
  assign n3095 = ~n2244 & n3094;
  assign n3096 = ~n1865 & ~n2242;
  assign n3097 = ~n3095 & n3096;
  assign n3098 = n1359 & n1368;
  assign n3099 = n2272 & n3098;
  assign n3100 = n2271 & n3099;
  assign n3101 = n2268 & n3100;
  assign n3102 = ~n1372 & n3101;
  assign n3103 = ~n2243 & n3102;
  assign n3104 = ~n2263 & n3103;
  assign n3105 = ~n966 & ~n1372;
  assign n3106 = ~n2243 & n3105;
  assign n3107 = ~n3104 & n3106;
  assign n3108 = ~pi087 & pi159;
  assign n3109 = pi087 & ~pi159;
  assign n3110 = ~pi088 & pi160;
  assign n3111 = pi088 & ~pi160;
  assign n3112 = ~pi089 & pi161;
  assign n3113 = pi089 & ~pi161;
  assign n3114 = ~pi090 & pi162;
  assign n3115 = pi090 & ~pi162;
  assign n3116 = ~pi091 & pi163;
  assign n3117 = pi091 & ~pi163;
  assign n3118 = ~pi092 & pi164;
  assign n3119 = pi092 & ~pi164;
  assign n3120 = pi094 & ~pi166;
  assign n3121 = pi093 & ~pi165;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = ~pi093 & pi165;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = ~n3119 & ~n3124;
  assign n3126 = ~n3118 & ~n3125;
  assign n3127 = ~n3117 & ~n3126;
  assign n3128 = ~n3116 & ~n3127;
  assign n3129 = ~n3115 & ~n3128;
  assign n3130 = ~n3114 & ~n3129;
  assign n3131 = ~n3113 & ~n3130;
  assign n3132 = ~n3112 & ~n3131;
  assign n3133 = ~n3111 & ~n3132;
  assign n3134 = ~n3110 & ~n3133;
  assign n3135 = ~n3109 & ~n3134;
  assign n3136 = ~n3108 & ~n3135;
  assign n3137 = ~pi087 & pi175;
  assign n3138 = pi087 & ~pi175;
  assign n3139 = ~pi088 & pi176;
  assign n3140 = pi088 & ~pi176;
  assign n3141 = ~pi089 & pi177;
  assign n3142 = pi089 & ~pi177;
  assign n3143 = ~pi090 & pi178;
  assign n3144 = pi090 & ~pi178;
  assign n3145 = ~pi091 & pi179;
  assign n3146 = pi091 & ~pi179;
  assign n3147 = ~pi092 & pi180;
  assign n3148 = pi092 & ~pi180;
  assign n3149 = pi094 & ~pi182;
  assign n3150 = pi093 & ~pi181;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = ~pi093 & pi181;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = ~n3148 & ~n3153;
  assign n3155 = ~n3147 & ~n3154;
  assign n3156 = ~n3146 & ~n3155;
  assign n3157 = ~n3145 & ~n3156;
  assign n3158 = ~n3144 & ~n3157;
  assign n3159 = ~n3143 & ~n3158;
  assign n3160 = ~n3142 & ~n3159;
  assign n3161 = ~n3141 & ~n3160;
  assign n3162 = ~n3140 & ~n3161;
  assign n3163 = ~n3139 & ~n3162;
  assign n3164 = ~n3138 & ~n3163;
  assign n3165 = ~n3137 & ~n3164;
  assign n3166 = ~n3136 & ~n3165;
  assign n3167 = ~pi087 & pi119;
  assign n3168 = pi087 & ~pi119;
  assign n3169 = ~pi088 & pi120;
  assign n3170 = pi088 & ~pi120;
  assign n3171 = ~pi089 & pi121;
  assign n3172 = pi089 & ~pi121;
  assign n3173 = ~pi090 & pi122;
  assign n3174 = pi090 & ~pi122;
  assign n3175 = ~pi091 & pi123;
  assign n3176 = pi091 & ~pi123;
  assign n3177 = ~pi092 & pi124;
  assign n3178 = pi092 & ~pi124;
  assign n3179 = pi094 & ~pi126;
  assign n3180 = pi093 & ~pi125;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~pi093 & pi125;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = ~n3178 & ~n3183;
  assign n3185 = ~n3177 & ~n3184;
  assign n3186 = ~n3176 & ~n3185;
  assign n3187 = ~n3175 & ~n3186;
  assign n3188 = ~n3174 & ~n3187;
  assign n3189 = ~n3173 & ~n3188;
  assign n3190 = ~n3172 & ~n3189;
  assign n3191 = ~n3171 & ~n3190;
  assign n3192 = ~n3170 & ~n3191;
  assign n3193 = ~n3169 & ~n3192;
  assign n3194 = ~n3168 & ~n3193;
  assign n3195 = ~n3167 & ~n3194;
  assign n3196 = ~pi087 & pi103;
  assign n3197 = pi087 & ~pi103;
  assign n3198 = ~pi088 & pi104;
  assign n3199 = pi088 & ~pi104;
  assign n3200 = ~pi089 & pi105;
  assign n3201 = pi089 & ~pi105;
  assign n3202 = ~pi090 & pi106;
  assign n3203 = pi090 & ~pi106;
  assign n3204 = ~pi091 & pi107;
  assign n3205 = pi091 & ~pi107;
  assign n3206 = ~pi092 & pi108;
  assign n3207 = pi092 & ~pi108;
  assign n3208 = pi094 & ~pi110;
  assign n3209 = pi093 & ~pi109;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = ~pi093 & pi109;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = ~n3207 & ~n3212;
  assign n3214 = ~n3206 & ~n3213;
  assign n3215 = ~n3205 & ~n3214;
  assign n3216 = ~n3204 & ~n3215;
  assign n3217 = ~n3203 & ~n3216;
  assign n3218 = ~n3202 & ~n3217;
  assign n3219 = ~n3201 & ~n3218;
  assign n3220 = ~n3200 & ~n3219;
  assign n3221 = ~n3199 & ~n3220;
  assign n3222 = ~n3198 & ~n3221;
  assign n3223 = ~n3197 & ~n3222;
  assign n3224 = ~n3196 & ~n3223;
  assign n3225 = ~n3195 & ~n3224;
  assign n3226 = n3166 & n3225;
  assign n3227 = ~pi087 & pi111;
  assign n3228 = pi089 & ~pi113;
  assign n3229 = ~pi090 & pi114;
  assign n3230 = pi090 & ~pi114;
  assign n3231 = ~pi091 & pi115;
  assign n3232 = pi091 & ~pi115;
  assign n3233 = ~pi092 & pi116;
  assign n3234 = pi092 & ~pi116;
  assign n3235 = pi094 & ~pi118;
  assign n3236 = pi093 & ~pi117;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = ~pi093 & pi117;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3234 & ~n3239;
  assign n3241 = ~n3233 & ~n3240;
  assign n3242 = ~n3232 & ~n3241;
  assign n3243 = ~n3231 & ~n3242;
  assign n3244 = ~n3230 & ~n3243;
  assign n3245 = ~n3229 & ~n3244;
  assign n3246 = ~n3228 & ~n3245;
  assign n3247 = ~pi089 & pi113;
  assign n3248 = ~pi088 & pi112;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n3246 & n3249;
  assign n3251 = pi087 & ~pi111;
  assign n3252 = pi088 & ~pi112;
  assign n3253 = ~n3251 & ~n3252;
  assign n3254 = ~n3250 & n3253;
  assign n3255 = ~n3227 & ~n3254;
  assign n3256 = ~pi087 & pi127;
  assign n3257 = pi089 & ~pi129;
  assign n3258 = ~pi090 & pi130;
  assign n3259 = pi090 & ~pi130;
  assign n3260 = ~pi091 & pi131;
  assign n3261 = pi091 & ~pi131;
  assign n3262 = ~pi092 & pi132;
  assign n3263 = pi092 & ~pi132;
  assign n3264 = pi094 & ~pi134;
  assign n3265 = pi093 & ~pi133;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~pi093 & pi133;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = ~n3263 & ~n3268;
  assign n3270 = ~n3262 & ~n3269;
  assign n3271 = ~n3261 & ~n3270;
  assign n3272 = ~n3260 & ~n3271;
  assign n3273 = ~n3259 & ~n3272;
  assign n3274 = ~n3258 & ~n3273;
  assign n3275 = ~n3257 & ~n3274;
  assign n3276 = ~pi089 & pi129;
  assign n3277 = ~pi088 & pi128;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n3275 & n3278;
  assign n3280 = pi087 & ~pi127;
  assign n3281 = pi088 & ~pi128;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = ~n3279 & n3282;
  assign n3284 = ~n3256 & ~n3283;
  assign n3285 = ~pi087 & pi095;
  assign n3286 = pi089 & ~pi097;
  assign n3287 = ~pi090 & pi098;
  assign n3288 = pi090 & ~pi098;
  assign n3289 = ~pi091 & pi099;
  assign n3290 = pi091 & ~pi099;
  assign n3291 = ~pi092 & pi100;
  assign n3292 = pi092 & ~pi100;
  assign n3293 = pi094 & ~pi102;
  assign n3294 = pi093 & ~pi101;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = ~pi093 & pi101;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n3292 & ~n3297;
  assign n3299 = ~n3291 & ~n3298;
  assign n3300 = ~n3290 & ~n3299;
  assign n3301 = ~n3289 & ~n3300;
  assign n3302 = ~n3288 & ~n3301;
  assign n3303 = ~n3287 & ~n3302;
  assign n3304 = ~n3286 & ~n3303;
  assign n3305 = ~pi089 & pi097;
  assign n3306 = ~pi088 & pi096;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = ~n3304 & n3307;
  assign n3309 = pi087 & ~pi095;
  assign n3310 = pi088 & ~pi096;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = ~n3308 & n3311;
  assign n3313 = ~n3285 & ~n3312;
  assign n3314 = ~n3284 & ~n3313;
  assign n3315 = ~n3255 & n3314;
  assign n3316 = ~pi087 & pi199;
  assign n3317 = pi089 & ~pi201;
  assign n3318 = ~pi090 & pi202;
  assign n3319 = pi090 & ~pi202;
  assign n3320 = ~pi091 & pi203;
  assign n3321 = pi091 & ~pi203;
  assign n3322 = ~pi092 & pi204;
  assign n3323 = pi092 & ~pi204;
  assign n3324 = pi094 & ~pi206;
  assign n3325 = pi093 & ~pi205;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = ~pi093 & pi205;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~n3323 & ~n3328;
  assign n3330 = ~n3322 & ~n3329;
  assign n3331 = ~n3321 & ~n3330;
  assign n3332 = ~n3320 & ~n3331;
  assign n3333 = ~n3319 & ~n3332;
  assign n3334 = ~n3318 & ~n3333;
  assign n3335 = ~n3317 & ~n3334;
  assign n3336 = ~pi089 & pi201;
  assign n3337 = ~pi088 & pi200;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = ~n3335 & n3338;
  assign n3340 = pi087 & ~pi199;
  assign n3341 = pi088 & ~pi200;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3339 & n3342;
  assign n3344 = ~n3316 & ~n3343;
  assign n3345 = ~pi087 & pi207;
  assign n3346 = pi089 & ~pi209;
  assign n3347 = ~pi090 & pi210;
  assign n3348 = pi090 & ~pi210;
  assign n3349 = ~pi091 & pi211;
  assign n3350 = pi091 & ~pi211;
  assign n3351 = ~pi092 & pi212;
  assign n3352 = pi092 & ~pi212;
  assign n3353 = pi094 & ~pi214;
  assign n3354 = pi093 & ~pi213;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = ~pi093 & pi213;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = ~n3352 & ~n3357;
  assign n3359 = ~n3351 & ~n3358;
  assign n3360 = ~n3350 & ~n3359;
  assign n3361 = ~n3349 & ~n3360;
  assign n3362 = ~n3348 & ~n3361;
  assign n3363 = ~n3347 & ~n3362;
  assign n3364 = ~n3346 & ~n3363;
  assign n3365 = ~pi089 & pi209;
  assign n3366 = ~pi088 & pi208;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = ~n3364 & n3367;
  assign n3369 = pi087 & ~pi207;
  assign n3370 = pi088 & ~pi208;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = ~n3368 & n3371;
  assign n3373 = ~n3345 & ~n3372;
  assign n3374 = ~n3344 & ~n3373;
  assign n3375 = ~pi087 & pi223;
  assign n3376 = pi089 & ~pi225;
  assign n3377 = ~pi090 & pi226;
  assign n3378 = pi090 & ~pi226;
  assign n3379 = ~pi091 & pi227;
  assign n3380 = pi091 & ~pi227;
  assign n3381 = ~pi092 & pi228;
  assign n3382 = pi092 & ~pi228;
  assign n3383 = pi094 & ~pi230;
  assign n3384 = pi093 & ~pi229;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = ~pi093 & pi229;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n3382 & ~n3387;
  assign n3389 = ~n3381 & ~n3388;
  assign n3390 = ~n3380 & ~n3389;
  assign n3391 = ~n3379 & ~n3390;
  assign n3392 = ~n3378 & ~n3391;
  assign n3393 = ~n3377 & ~n3392;
  assign n3394 = ~n3376 & ~n3393;
  assign n3395 = ~pi089 & pi225;
  assign n3396 = ~pi088 & pi224;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3394 & n3397;
  assign n3399 = pi087 & ~pi223;
  assign n3400 = pi088 & ~pi224;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~n3398 & n3401;
  assign n3403 = ~n3375 & ~n3402;
  assign n3404 = ~pi087 & pi151;
  assign n3405 = pi089 & ~pi153;
  assign n3406 = ~pi090 & pi154;
  assign n3407 = pi090 & ~pi154;
  assign n3408 = ~pi091 & pi155;
  assign n3409 = pi091 & ~pi155;
  assign n3410 = ~pi092 & pi156;
  assign n3411 = pi092 & ~pi156;
  assign n3412 = pi094 & ~pi158;
  assign n3413 = pi093 & ~pi157;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~pi093 & pi157;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~n3411 & ~n3416;
  assign n3418 = ~n3410 & ~n3417;
  assign n3419 = ~n3409 & ~n3418;
  assign n3420 = ~n3408 & ~n3419;
  assign n3421 = ~n3407 & ~n3420;
  assign n3422 = ~n3406 & ~n3421;
  assign n3423 = ~n3405 & ~n3422;
  assign n3424 = ~pi089 & pi153;
  assign n3425 = ~pi088 & pi152;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = ~n3423 & n3426;
  assign n3428 = pi087 & ~pi151;
  assign n3429 = pi088 & ~pi152;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = ~n3427 & n3430;
  assign n3432 = ~n3404 & ~n3431;
  assign n3433 = ~n3403 & ~n3432;
  assign n3434 = n3374 & n3433;
  assign n3435 = n3315 & n3434;
  assign n3436 = ~pi087 & pi191;
  assign n3437 = pi087 & ~pi191;
  assign n3438 = ~pi088 & pi192;
  assign n3439 = pi088 & ~pi192;
  assign n3440 = ~pi089 & pi193;
  assign n3441 = pi089 & ~pi193;
  assign n3442 = ~pi090 & pi194;
  assign n3443 = pi090 & ~pi194;
  assign n3444 = ~pi091 & pi195;
  assign n3445 = pi091 & ~pi195;
  assign n3446 = ~pi092 & pi196;
  assign n3447 = pi092 & ~pi196;
  assign n3448 = pi094 & ~pi198;
  assign n3449 = pi093 & ~pi197;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~pi093 & pi197;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = ~n3447 & ~n3452;
  assign n3454 = ~n3446 & ~n3453;
  assign n3455 = ~n3445 & ~n3454;
  assign n3456 = ~n3444 & ~n3455;
  assign n3457 = ~n3443 & ~n3456;
  assign n3458 = ~n3442 & ~n3457;
  assign n3459 = ~n3441 & ~n3458;
  assign n3460 = ~n3440 & ~n3459;
  assign n3461 = ~n3439 & ~n3460;
  assign n3462 = ~n3438 & ~n3461;
  assign n3463 = ~n3437 & ~n3462;
  assign n3464 = ~n3436 & ~n3463;
  assign n3465 = ~pi087 & pi143;
  assign n3466 = pi087 & ~pi143;
  assign n3467 = ~pi088 & pi144;
  assign n3468 = pi088 & ~pi144;
  assign n3469 = ~pi089 & pi145;
  assign n3470 = pi089 & ~pi145;
  assign n3471 = ~pi090 & pi146;
  assign n3472 = pi090 & ~pi146;
  assign n3473 = ~pi091 & pi147;
  assign n3474 = pi091 & ~pi147;
  assign n3475 = ~pi092 & pi148;
  assign n3476 = pi092 & ~pi148;
  assign n3477 = pi094 & ~pi150;
  assign n3478 = pi093 & ~pi149;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = ~pi093 & pi149;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = ~n3476 & ~n3481;
  assign n3483 = ~n3475 & ~n3482;
  assign n3484 = ~n3474 & ~n3483;
  assign n3485 = ~n3473 & ~n3484;
  assign n3486 = ~n3472 & ~n3485;
  assign n3487 = ~n3471 & ~n3486;
  assign n3488 = ~n3470 & ~n3487;
  assign n3489 = ~n3469 & ~n3488;
  assign n3490 = ~n3468 & ~n3489;
  assign n3491 = ~n3467 & ~n3490;
  assign n3492 = ~n3466 & ~n3491;
  assign n3493 = ~n3465 & ~n3492;
  assign n3494 = ~n3464 & ~n3493;
  assign n3495 = n3435 & n3494;
  assign n3496 = ~pi087 & pi183;
  assign n3497 = pi089 & ~pi185;
  assign n3498 = ~pi090 & pi186;
  assign n3499 = pi090 & ~pi186;
  assign n3500 = ~pi091 & pi187;
  assign n3501 = pi091 & ~pi187;
  assign n3502 = ~pi092 & pi188;
  assign n3503 = pi092 & ~pi188;
  assign n3504 = pi094 & ~pi190;
  assign n3505 = pi093 & ~pi189;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = ~pi093 & pi189;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3503 & ~n3508;
  assign n3510 = ~n3502 & ~n3509;
  assign n3511 = ~n3501 & ~n3510;
  assign n3512 = ~n3500 & ~n3511;
  assign n3513 = ~n3499 & ~n3512;
  assign n3514 = ~n3498 & ~n3513;
  assign n3515 = ~n3497 & ~n3514;
  assign n3516 = ~pi089 & pi185;
  assign n3517 = ~pi088 & pi184;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~n3515 & n3518;
  assign n3520 = pi087 & ~pi183;
  assign n3521 = pi088 & ~pi184;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = ~n3519 & n3522;
  assign n3524 = ~n3496 & ~n3523;
  assign n3525 = ~pi087 & pi135;
  assign n3526 = pi089 & ~pi137;
  assign n3527 = ~pi090 & pi138;
  assign n3528 = pi090 & ~pi138;
  assign n3529 = ~pi091 & pi139;
  assign n3530 = pi091 & ~pi139;
  assign n3531 = ~pi092 & pi140;
  assign n3532 = pi092 & ~pi140;
  assign n3533 = pi094 & ~pi142;
  assign n3534 = pi093 & ~pi141;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~pi093 & pi141;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n3532 & ~n3537;
  assign n3539 = ~n3531 & ~n3538;
  assign n3540 = ~n3530 & ~n3539;
  assign n3541 = ~n3529 & ~n3540;
  assign n3542 = ~n3528 & ~n3541;
  assign n3543 = ~n3527 & ~n3542;
  assign n3544 = ~n3526 & ~n3543;
  assign n3545 = ~pi089 & pi137;
  assign n3546 = ~pi088 & pi136;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = ~n3544 & n3547;
  assign n3549 = pi087 & ~pi135;
  assign n3550 = pi088 & ~pi136;
  assign n3551 = ~n3549 & ~n3550;
  assign n3552 = ~n3548 & n3551;
  assign n3553 = ~n3525 & ~n3552;
  assign n3554 = ~n3524 & ~n3553;
  assign n3555 = n2317 & n3554;
  assign n3556 = pi007 & ~n501;
  assign n3557 = n2311 & n3556;
  assign n3558 = n2309 & n3557;
  assign n3559 = ~n2306 & n3558;
  assign n3560 = ~n500 & n3559;
  assign n3561 = n2316 & n3560;
  assign n3562 = n3555 & n3561;
  assign n3563 = ~pi087 & pi255;
  assign n3564 = pi089 & ~pi257;
  assign n3565 = ~pi090 & pi258;
  assign n3566 = pi090 & ~pi258;
  assign n3567 = ~pi091 & pi259;
  assign n3568 = pi091 & ~pi259;
  assign n3569 = ~pi092 & pi260;
  assign n3570 = pi092 & ~pi260;
  assign n3571 = pi094 & ~pi262;
  assign n3572 = pi093 & ~pi261;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = ~pi093 & pi261;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = ~n3570 & ~n3575;
  assign n3577 = ~n3569 & ~n3576;
  assign n3578 = ~n3568 & ~n3577;
  assign n3579 = ~n3567 & ~n3578;
  assign n3580 = ~n3566 & ~n3579;
  assign n3581 = ~n3565 & ~n3580;
  assign n3582 = ~n3564 & ~n3581;
  assign n3583 = ~pi089 & pi257;
  assign n3584 = ~pi088 & pi256;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = ~n3582 & n3585;
  assign n3587 = pi087 & ~pi255;
  assign n3588 = pi088 & ~pi256;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3586 & n3589;
  assign n3591 = ~n3563 & ~n3590;
  assign n3592 = ~pi087 & pi247;
  assign n3593 = pi089 & ~pi249;
  assign n3594 = ~pi090 & pi250;
  assign n3595 = pi090 & ~pi250;
  assign n3596 = ~pi091 & pi251;
  assign n3597 = pi091 & ~pi251;
  assign n3598 = ~pi092 & pi252;
  assign n3599 = pi092 & ~pi252;
  assign n3600 = pi094 & ~pi254;
  assign n3601 = pi093 & ~pi253;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = ~pi093 & pi253;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = ~n3599 & ~n3604;
  assign n3606 = ~n3598 & ~n3605;
  assign n3607 = ~n3597 & ~n3606;
  assign n3608 = ~n3596 & ~n3607;
  assign n3609 = ~n3595 & ~n3608;
  assign n3610 = ~n3594 & ~n3609;
  assign n3611 = ~n3593 & ~n3610;
  assign n3612 = ~pi089 & pi249;
  assign n3613 = ~pi088 & pi248;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = ~n3611 & n3614;
  assign n3616 = pi087 & ~pi247;
  assign n3617 = pi088 & ~pi248;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = ~n3615 & n3618;
  assign n3620 = ~n3592 & ~n3619;
  assign n3621 = ~n3591 & ~n3620;
  assign n3622 = ~pi087 & pi263;
  assign n3623 = pi089 & ~pi265;
  assign n3624 = ~pi090 & pi266;
  assign n3625 = pi090 & ~pi266;
  assign n3626 = ~pi091 & pi267;
  assign n3627 = pi091 & ~pi267;
  assign n3628 = ~pi092 & pi268;
  assign n3629 = pi092 & ~pi268;
  assign n3630 = pi094 & ~pi270;
  assign n3631 = pi093 & ~pi269;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = ~pi093 & pi269;
  assign n3634 = ~n3632 & ~n3633;
  assign n3635 = ~n3629 & ~n3634;
  assign n3636 = ~n3628 & ~n3635;
  assign n3637 = ~n3627 & ~n3636;
  assign n3638 = ~n3626 & ~n3637;
  assign n3639 = ~n3625 & ~n3638;
  assign n3640 = ~n3624 & ~n3639;
  assign n3641 = ~n3623 & ~n3640;
  assign n3642 = ~pi089 & pi265;
  assign n3643 = ~pi088 & pi264;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = ~n3641 & n3644;
  assign n3646 = pi087 & ~pi263;
  assign n3647 = pi088 & ~pi264;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = ~n3645 & n3648;
  assign n3650 = ~n3622 & ~n3649;
  assign n3651 = ~pi087 & pi167;
  assign n3652 = pi089 & ~pi169;
  assign n3653 = ~pi090 & pi170;
  assign n3654 = pi090 & ~pi170;
  assign n3655 = ~pi091 & pi171;
  assign n3656 = pi091 & ~pi171;
  assign n3657 = ~pi092 & pi172;
  assign n3658 = pi092 & ~pi172;
  assign n3659 = pi094 & ~pi174;
  assign n3660 = pi093 & ~pi173;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = ~pi093 & pi173;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = ~n3658 & ~n3663;
  assign n3665 = ~n3657 & ~n3664;
  assign n3666 = ~n3656 & ~n3665;
  assign n3667 = ~n3655 & ~n3666;
  assign n3668 = ~n3654 & ~n3667;
  assign n3669 = ~n3653 & ~n3668;
  assign n3670 = ~n3652 & ~n3669;
  assign n3671 = ~pi089 & pi169;
  assign n3672 = ~pi088 & pi168;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = ~n3670 & n3673;
  assign n3675 = pi087 & ~pi167;
  assign n3676 = pi088 & ~pi168;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3674 & n3677;
  assign n3679 = ~n3651 & ~n3678;
  assign n3680 = ~n3650 & ~n3679;
  assign n3681 = n3621 & n3680;
  assign n3682 = ~pi087 & pi271;
  assign n3683 = pi089 & ~pi273;
  assign n3684 = ~pi090 & pi274;
  assign n3685 = pi090 & ~pi274;
  assign n3686 = ~pi091 & pi275;
  assign n3687 = pi091 & ~pi275;
  assign n3688 = ~pi092 & pi276;
  assign n3689 = pi092 & ~pi276;
  assign n3690 = pi094 & ~pi278;
  assign n3691 = pi093 & ~pi277;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = ~pi093 & pi277;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~n3689 & ~n3694;
  assign n3696 = ~n3688 & ~n3695;
  assign n3697 = ~n3687 & ~n3696;
  assign n3698 = ~n3686 & ~n3697;
  assign n3699 = ~n3685 & ~n3698;
  assign n3700 = ~n3684 & ~n3699;
  assign n3701 = ~n3683 & ~n3700;
  assign n3702 = ~pi089 & pi273;
  assign n3703 = ~pi088 & pi272;
  assign n3704 = ~n3702 & ~n3703;
  assign n3705 = ~n3701 & n3704;
  assign n3706 = pi087 & ~pi271;
  assign n3707 = pi088 & ~pi272;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = ~n3705 & n3708;
  assign n3710 = ~n3682 & ~n3709;
  assign n3711 = ~pi087 & pi239;
  assign n3712 = pi089 & ~pi241;
  assign n3713 = ~pi090 & pi242;
  assign n3714 = pi090 & ~pi242;
  assign n3715 = ~pi091 & pi243;
  assign n3716 = pi091 & ~pi243;
  assign n3717 = ~pi092 & pi244;
  assign n3718 = pi092 & ~pi244;
  assign n3719 = pi094 & ~pi246;
  assign n3720 = pi093 & ~pi245;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = ~pi093 & pi245;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3718 & ~n3723;
  assign n3725 = ~n3717 & ~n3724;
  assign n3726 = ~n3716 & ~n3725;
  assign n3727 = ~n3715 & ~n3726;
  assign n3728 = ~n3714 & ~n3727;
  assign n3729 = ~n3713 & ~n3728;
  assign n3730 = ~n3712 & ~n3729;
  assign n3731 = ~pi089 & pi241;
  assign n3732 = ~pi088 & pi240;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n3730 & n3733;
  assign n3735 = pi087 & ~pi239;
  assign n3736 = pi088 & ~pi240;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = ~n3734 & n3737;
  assign n3739 = ~n3711 & ~n3738;
  assign n3740 = ~n3710 & ~n3739;
  assign n3741 = ~pi087 & pi231;
  assign n3742 = pi089 & ~pi233;
  assign n3743 = ~pi090 & pi234;
  assign n3744 = pi090 & ~pi234;
  assign n3745 = ~pi091 & pi235;
  assign n3746 = pi091 & ~pi235;
  assign n3747 = ~pi092 & pi236;
  assign n3748 = pi092 & ~pi236;
  assign n3749 = pi094 & ~pi238;
  assign n3750 = pi093 & ~pi237;
  assign n3751 = ~n3749 & ~n3750;
  assign n3752 = ~pi093 & pi237;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = ~n3748 & ~n3753;
  assign n3755 = ~n3747 & ~n3754;
  assign n3756 = ~n3746 & ~n3755;
  assign n3757 = ~n3745 & ~n3756;
  assign n3758 = ~n3744 & ~n3757;
  assign n3759 = ~n3743 & ~n3758;
  assign n3760 = ~n3742 & ~n3759;
  assign n3761 = ~pi089 & pi233;
  assign n3762 = ~pi088 & pi232;
  assign n3763 = ~n3761 & ~n3762;
  assign n3764 = ~n3760 & n3763;
  assign n3765 = pi087 & ~pi231;
  assign n3766 = pi088 & ~pi232;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = ~n3764 & n3767;
  assign n3769 = ~n3741 & ~n3768;
  assign n3770 = ~pi087 & pi215;
  assign n3771 = pi089 & ~pi217;
  assign n3772 = ~pi090 & pi218;
  assign n3773 = pi090 & ~pi218;
  assign n3774 = ~pi091 & pi219;
  assign n3775 = pi091 & ~pi219;
  assign n3776 = ~pi092 & pi220;
  assign n3777 = pi092 & ~pi220;
  assign n3778 = pi094 & ~pi222;
  assign n3779 = pi093 & ~pi221;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = ~pi093 & pi221;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~n3777 & ~n3782;
  assign n3784 = ~n3776 & ~n3783;
  assign n3785 = ~n3775 & ~n3784;
  assign n3786 = ~n3774 & ~n3785;
  assign n3787 = ~n3773 & ~n3786;
  assign n3788 = ~n3772 & ~n3787;
  assign n3789 = ~n3771 & ~n3788;
  assign n3790 = ~pi089 & pi217;
  assign n3791 = ~pi088 & pi216;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = ~n3789 & n3792;
  assign n3794 = pi087 & ~pi215;
  assign n3795 = pi088 & ~pi216;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = ~n3793 & n3796;
  assign n3798 = ~n3770 & ~n3797;
  assign n3799 = ~n3769 & ~n3798;
  assign n3800 = n3740 & n3799;
  assign n3801 = n3681 & n3800;
  assign n3802 = n3562 & n3801;
  assign n3803 = n3495 & n3802;
  assign n3804 = n3226 & n3803;
  assign n3805 = ~n3107 & n3804;
  assign n3806 = ~n3097 & n3805;
  assign n3807 = ~n3067 & n3806;
  assign n3808 = ~n1463 & ~n2110;
  assign n3809 = ~n1493 & n3808;
  assign n3810 = ~n2307 & ~n2364;
  assign n3811 = ~n3285 & n3810;
  assign n3812 = ~n534 & ~n2082;
  assign n3813 = n2308 & n3812;
  assign n3814 = pi008 & ~n501;
  assign n3815 = n2311 & n3814;
  assign n3816 = n3813 & n3815;
  assign n3817 = n3811 & n3816;
  assign n3818 = ~n2306 & n3817;
  assign n3819 = ~n2391 & ~n3312;
  assign n3820 = n3818 & n3819;
  assign n3821 = ~n500 & ~n532;
  assign n3822 = ~n562 & ~n594;
  assign n3823 = n3821 & n3822;
  assign n3824 = n3820 & n3823;
  assign n3825 = n3809 & n3824;
  assign n3826 = ~n2245 & ~po145;
  assign n3827 = ~n2324 & n3826;
  assign n3828 = ~n2322 & n3827;
  assign n3829 = n2325 & ~n3828;
  assign n3830 = ~n2242 & ~n3095;
  assign n3831 = ~n1372 & ~n2243;
  assign n3832 = ~n3104 & n3831;
  assign n3833 = ~n3830 & ~n3832;
  assign n3834 = n3829 & n3833;
  assign n3835 = ~n3825 & ~n3834;
  assign n3836 = ~n3807 & n3835;
  assign n3837 = ~po145 & ~n3828;
  assign n3838 = ~n2663 & ~n2842;
  assign n3839 = ~n2692 & ~n2722;
  assign n3840 = n3838 & n3839;
  assign n3841 = ~n2965 & n3840;
  assign n3842 = ~n2994 & ~n3024;
  assign n3843 = n3841 & n3842;
  assign n3844 = pi005 & ~n2363;
  assign n3845 = ~n2392 & ~n2543;
  assign n3846 = ~n2572 & ~n2602;
  assign n3847 = n3845 & n3846;
  assign n3848 = n3844 & n3847;
  assign n3849 = ~n2512 & ~n2754;
  assign n3850 = ~n2783 & ~n2813;
  assign n3851 = n3849 & n3850;
  assign n3852 = ~n2424 & ~n2631;
  assign n3853 = ~n2453 & ~n2483;
  assign n3854 = n3852 & n3853;
  assign n3855 = n3851 & n3854;
  assign n3856 = n3848 & n3855;
  assign n3857 = n3843 & n3856;
  assign n3858 = ~n504 & ~n1435;
  assign n3859 = ~n1465 & ~n2307;
  assign n3860 = n3858 & n3859;
  assign n3861 = n2246 & n3860;
  assign n3862 = ~n2306 & n3861;
  assign n3863 = ~n500 & n3862;
  assign n3864 = n2318 & n3863;
  assign n3865 = n2723 & ~n3864;
  assign n3866 = ~n2905 & ~n3053;
  assign n3867 = ~n2876 & ~n2934;
  assign n3868 = n3866 & n3867;
  assign n3869 = ~n3865 & n3868;
  assign n3870 = n3857 & n3869;
  assign n3871 = ~n3066 & n3870;
  assign n3872 = n2331 & ~n3104;
  assign n3873 = n2329 & ~n3095;
  assign n3874 = ~n3872 & ~n3873;
  assign n3875 = n3871 & n3874;
  assign n3876 = ~n3837 & n3875;
  assign n3877 = n1774 & ~n3065;
  assign n3878 = n2244 & ~n3104;
  assign n3879 = n1680 & n2112;
  assign n3880 = n2051 & n2207;
  assign n3881 = n3879 & n3880;
  assign n3882 = n1434 & n1618;
  assign n3883 = n1557 & n1741;
  assign n3884 = n3882 & n3883;
  assign n3885 = n3881 & n3884;
  assign n3886 = n1464 & ~n3864;
  assign n3887 = ~n1804 & ~n1988;
  assign n3888 = n1866 & n3887;
  assign n3889 = ~n1897 & n2254;
  assign n3890 = n3082 & n3889;
  assign n3891 = n3888 & n3890;
  assign n3892 = ~n3886 & n3891;
  assign n3893 = n3885 & n3892;
  assign n3894 = ~n2242 & n3893;
  assign n3895 = ~n3095 & n3894;
  assign n3896 = ~n3878 & n3895;
  assign n3897 = ~n3877 & n3896;
  assign n3898 = ~n3837 & n3897;
  assign n3899 = ~n3876 & ~n3898;
  assign n3900 = n905 & ~n3066;
  assign n3901 = n2263 & ~n3094;
  assign n3902 = ~n563 & n719;
  assign n3903 = n2266 & n3902;
  assign n3904 = n2274 & n3903;
  assign n3905 = n533 & ~n3864;
  assign n3906 = ~n966 & n2269;
  assign n3907 = ~n3905 & n3906;
  assign n3908 = n3904 & n3907;
  assign n3909 = ~n1372 & n3908;
  assign n3910 = ~n2243 & n3909;
  assign n3911 = ~n3104 & n3910;
  assign n3912 = ~n3901 & n3911;
  assign n3913 = ~n3837 & n3912;
  assign n3914 = ~n3900 & n3913;
  assign n3915 = ~n1464 & ~n2242;
  assign n3916 = ~n3095 & n3915;
  assign n3917 = ~n533 & ~n1372;
  assign n3918 = ~n2243 & n3917;
  assign n3919 = ~n3104 & n3918;
  assign n3920 = pi006 & ~n3864;
  assign n3921 = ~n3919 & n3920;
  assign n3922 = ~n3916 & n3921;
  assign n3923 = ~n2723 & ~n3066;
  assign n3924 = ~n3837 & ~n3923;
  assign n3925 = n3922 & n3924;
  assign n3926 = ~n3914 & ~n3925;
  assign n3927 = n3899 & n3926;
  assign po004 = ~n3836 | ~n3927;
  assign n3929 = ~n3864 & ~n3919;
  assign n3930 = ~n3916 & n3929;
  assign n3931 = n3924 & n3930;
  assign n3932 = ~n3864 & ~n3931;
  assign n3933 = n2316 & n3863;
  assign n3934 = n3555 & n3933;
  assign n3935 = n3801 & n3934;
  assign n3936 = n3495 & n3935;
  assign n3937 = n3226 & n3936;
  assign n3938 = ~n3107 & n3937;
  assign n3939 = ~n3097 & n3938;
  assign n3940 = ~n3067 & n3939;
  assign n3941 = ~n2364 & ~n3285;
  assign n3942 = n3859 & n3941;
  assign n3943 = n3812 & n3858;
  assign n3944 = n2246 & n3943;
  assign n3945 = n3942 & n3944;
  assign n3946 = ~n2306 & n3945;
  assign n3947 = n3819 & n3946;
  assign n3948 = n3823 & n3947;
  assign po149 = n3809 & n3948;
  assign n3950 = n3313 & ~po149;
  assign n3951 = n3621 & n3799;
  assign n3952 = n3554 & n3740;
  assign n3953 = n3951 & n3952;
  assign n3954 = ~n3255 & ~n3284;
  assign n3955 = n3433 & n3954;
  assign n3956 = n3374 & n3680;
  assign n3957 = n3955 & n3956;
  assign n3958 = n3494 & n3957;
  assign n3959 = n3953 & n3958;
  assign n3960 = n3226 & n3959;
  assign n3961 = ~n3950 & n3960;
  assign n3962 = ~n3940 & n3961;
  assign n3963 = ~n3932 & n3962;
  assign n3964 = n3099 & n3903;
  assign n3965 = n3907 & n3964;
  assign n3966 = ~n1372 & n3965;
  assign n3967 = ~n2243 & n3966;
  assign n3968 = ~n3104 & n3967;
  assign n3969 = ~n3901 & n3968;
  assign n3970 = ~n3837 & n3969;
  assign n3971 = ~n3900 & n3970;
  assign n3972 = n3107 & ~n3971;
  assign n3973 = n2693 & ~n2722;
  assign n3974 = ~n2965 & n3973;
  assign n3975 = n3842 & n3974;
  assign n3976 = n2393 & n2633;
  assign n3977 = n2514 & n2844;
  assign n3978 = n3976 & n3977;
  assign n3979 = n3975 & n3978;
  assign n3980 = n3869 & n3979;
  assign n3981 = ~n3066 & n3980;
  assign n3982 = n3874 & n3981;
  assign n3983 = ~n3837 & n3982;
  assign n3984 = n3067 & ~n3983;
  assign n3985 = n3073 & n3087;
  assign n3986 = ~n1433 & n3075;
  assign n3987 = n3070 & n3986;
  assign n3988 = n3985 & n3987;
  assign n3989 = n3082 & n3089;
  assign n3990 = n3888 & n3989;
  assign n3991 = ~n3886 & n3990;
  assign n3992 = n3988 & n3991;
  assign n3993 = ~n2242 & n3992;
  assign n3994 = ~n3095 & n3993;
  assign n3995 = ~n3878 & n3994;
  assign n3996 = ~n3877 & n3995;
  assign n3997 = ~n3837 & n3996;
  assign n3998 = n3097 & ~n3997;
  assign n3999 = ~n3984 & ~n3998;
  assign n4000 = ~n3972 & n3999;
  assign n4001 = n3963 & n4000;
  assign n4002 = n3833 & n3837;
  assign n4003 = n3837 & ~n4002;
  assign n4004 = n2392 & ~po149;
  assign n4005 = ~n2363 & ~n2543;
  assign n4006 = n3846 & n4005;
  assign n4007 = n3854 & n4006;
  assign n4008 = n3840 & n3851;
  assign n4009 = ~n2965 & ~n3024;
  assign n4010 = n4008 & n4009;
  assign n4011 = n4007 & n4010;
  assign n4012 = n3868 & n4011;
  assign n4013 = ~n4004 & n4012;
  assign n4014 = ~n3066 & n4013;
  assign n4015 = ~n3983 & n4014;
  assign n4016 = ~n4003 & n4015;
  assign n4017 = n3873 & ~n3997;
  assign n4018 = n2994 & ~n3940;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = n3872 & ~n3971;
  assign n4021 = n3865 & ~n3931;
  assign n4022 = ~n4020 & ~n4021;
  assign n4023 = n4019 & n4022;
  assign n4024 = n4016 & n4023;
  assign n4025 = n2111 & ~po149;
  assign n4026 = ~n1649 & ~n2081;
  assign n4027 = n3072 & n4026;
  assign n4028 = n3880 & n4027;
  assign n4029 = n3987 & n4028;
  assign n4030 = ~n1835 & n3887;
  assign n4031 = n3890 & n4030;
  assign n4032 = n4029 & n4031;
  assign n4033 = ~n4025 & n4032;
  assign n4034 = ~n2242 & n4033;
  assign n4035 = ~n3095 & n4034;
  assign n4036 = ~n3997 & n4035;
  assign n4037 = ~n4003 & n4036;
  assign n4038 = n3877 & ~n3983;
  assign n4039 = n3878 & ~n3971;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = n1865 & ~n3940;
  assign n4042 = n3886 & ~n3931;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = n4040 & n4043;
  assign n4045 = n4037 & n4044;
  assign n4046 = n3901 & ~n3997;
  assign n4047 = n563 & ~po149;
  assign n4048 = ~n875 & n1360;
  assign n4049 = n843 & n1240;
  assign n4050 = n720 & n4049;
  assign n4051 = n4048 & n4050;
  assign n4052 = ~n4047 & n4051;
  assign n4053 = n3831 & n4052;
  assign n4054 = ~n3104 & n4053;
  assign n4055 = ~n3837 & n4054;
  assign n4056 = ~n3971 & n4055;
  assign n4057 = ~n4046 & n4056;
  assign n4058 = n3905 & ~n3931;
  assign n4059 = n3900 & ~n3983;
  assign n4060 = n966 & ~n3940;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = ~n4058 & n4061;
  assign n4063 = n4057 & n4062;
  assign n4064 = ~n4045 & ~n4063;
  assign n4065 = ~n4024 & ~n4064;
  assign n4066 = n3920 & ~n3931;
  assign n4067 = ~n4003 & n4066;
  assign n4068 = n3923 & ~n3983;
  assign n4069 = n3919 & ~n3971;
  assign n4070 = n3916 & ~n3997;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = ~n4068 & n4071;
  assign n4073 = n4067 & n4072;
  assign n4074 = n3054 & n3974;
  assign n4075 = n2633 & n3844;
  assign n4076 = n3977 & n4075;
  assign n4077 = n4074 & n4076;
  assign n4078 = n2936 & n4077;
  assign n4079 = ~n4004 & n4078;
  assign n4080 = ~n3066 & n4079;
  assign n4081 = ~n3983 & n4080;
  assign n4082 = ~n4003 & n4081;
  assign n4083 = n4023 & n4082;
  assign n4084 = ~n4073 & ~n4083;
  assign n4085 = ~n4065 & n4084;
  assign n4086 = ~n4001 & ~n4085;
  assign n4087 = ~n3165 & ~n3195;
  assign n4088 = ~n3224 & n4087;
  assign n4089 = ~n3284 & ~n3432;
  assign n4090 = ~n3255 & n4089;
  assign n4091 = ~n3464 & n4090;
  assign n4092 = ~n3136 & ~n3493;
  assign n4093 = n4091 & n4092;
  assign n4094 = pi007 & ~n3524;
  assign n4095 = ~n3553 & ~n3710;
  assign n4096 = ~n3739 & ~n3769;
  assign n4097 = n4095 & n4096;
  assign n4098 = n4094 & n4097;
  assign n4099 = ~n3344 & ~n3679;
  assign n4100 = ~n3373 & ~n3403;
  assign n4101 = n4099 & n4100;
  assign n4102 = ~n3591 & ~n3798;
  assign n4103 = ~n3620 & ~n3650;
  assign n4104 = n4102 & n4103;
  assign n4105 = n4101 & n4104;
  assign n4106 = n4098 & n4105;
  assign n4107 = n4093 & n4106;
  assign n4108 = n4088 & n4107;
  assign n4109 = ~n3950 & n4108;
  assign n4110 = ~n3940 & n4109;
  assign n4111 = ~n3932 & n4110;
  assign n4112 = n4000 & n4111;
  assign n4113 = ~n4086 & ~n4112;
  assign n4114 = ~n3932 & ~po149;
  assign n4115 = ~n2392 & ~n3066;
  assign n4116 = ~n3983 & n4115;
  assign n4117 = ~n2111 & ~n2242;
  assign n4118 = ~n3095 & n4117;
  assign n4119 = ~n3997 & n4118;
  assign n4120 = ~n4116 & ~n4119;
  assign n4121 = ~n563 & ~n1372;
  assign n4122 = ~n2243 & n4121;
  assign n4123 = ~n3104 & n4122;
  assign n4124 = ~n3971 & n4123;
  assign n4125 = ~n3313 & ~n3940;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = n4120 & n4126;
  assign n4128 = n4114 & n4127;
  assign n4129 = ~n4113 & ~n4128;
  assign n4130 = pi008 & ~po149;
  assign n4131 = ~n3932 & n4130;
  assign n4132 = n4127 & n4131;
  assign n4133 = ~n2905 & ~n3066;
  assign n4134 = ~n3983 & n4133;
  assign n4135 = ~pi103 & pi175;
  assign n4136 = pi103 & ~pi175;
  assign n4137 = ~pi104 & pi176;
  assign n4138 = pi104 & ~pi176;
  assign n4139 = ~pi105 & pi177;
  assign n4140 = pi105 & ~pi177;
  assign n4141 = ~pi106 & pi178;
  assign n4142 = pi106 & ~pi178;
  assign n4143 = ~pi107 & pi179;
  assign n4144 = pi107 & ~pi179;
  assign n4145 = ~pi108 & pi180;
  assign n4146 = pi108 & ~pi180;
  assign n4147 = pi110 & ~pi182;
  assign n4148 = pi109 & ~pi181;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = ~pi109 & pi181;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = ~n4146 & ~n4151;
  assign n4153 = ~n4145 & ~n4152;
  assign n4154 = ~n4144 & ~n4153;
  assign n4155 = ~n4143 & ~n4154;
  assign n4156 = ~n4142 & ~n4155;
  assign n4157 = ~n4141 & ~n4156;
  assign n4158 = ~n4140 & ~n4157;
  assign n4159 = ~n4139 & ~n4158;
  assign n4160 = ~n4138 & ~n4159;
  assign n4161 = ~n4137 & ~n4160;
  assign n4162 = ~n4136 & ~n4161;
  assign n4163 = ~n4135 & ~n4162;
  assign n4164 = ~pi103 & pi191;
  assign n4165 = pi103 & ~pi191;
  assign n4166 = ~pi104 & pi192;
  assign n4167 = pi104 & ~pi192;
  assign n4168 = ~pi105 & pi193;
  assign n4169 = pi105 & ~pi193;
  assign n4170 = ~pi106 & pi194;
  assign n4171 = pi106 & ~pi194;
  assign n4172 = ~pi107 & pi195;
  assign n4173 = pi107 & ~pi195;
  assign n4174 = ~pi108 & pi196;
  assign n4175 = pi108 & ~pi196;
  assign n4176 = pi110 & ~pi198;
  assign n4177 = pi109 & ~pi197;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = ~pi109 & pi197;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = ~n4175 & ~n4180;
  assign n4182 = ~n4174 & ~n4181;
  assign n4183 = ~n4173 & ~n4182;
  assign n4184 = ~n4172 & ~n4183;
  assign n4185 = ~n4171 & ~n4184;
  assign n4186 = ~n4170 & ~n4185;
  assign n4187 = ~n4169 & ~n4186;
  assign n4188 = ~n4168 & ~n4187;
  assign n4189 = ~n4167 & ~n4188;
  assign n4190 = ~n4166 & ~n4189;
  assign n4191 = ~n4165 & ~n4190;
  assign n4192 = ~n4164 & ~n4191;
  assign n4193 = ~n4163 & ~n4192;
  assign n4194 = ~pi103 & pi143;
  assign n4195 = pi103 & ~pi143;
  assign n4196 = ~pi104 & pi144;
  assign n4197 = pi104 & ~pi144;
  assign n4198 = ~pi105 & pi145;
  assign n4199 = pi105 & ~pi145;
  assign n4200 = ~pi106 & pi146;
  assign n4201 = pi106 & ~pi146;
  assign n4202 = ~pi107 & pi147;
  assign n4203 = pi107 & ~pi147;
  assign n4204 = ~pi108 & pi148;
  assign n4205 = pi108 & ~pi148;
  assign n4206 = pi110 & ~pi150;
  assign n4207 = pi109 & ~pi149;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = ~pi109 & pi149;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = ~n4205 & ~n4210;
  assign n4212 = ~n4204 & ~n4211;
  assign n4213 = ~n4203 & ~n4212;
  assign n4214 = ~n4202 & ~n4213;
  assign n4215 = ~n4201 & ~n4214;
  assign n4216 = ~n4200 & ~n4215;
  assign n4217 = ~n4199 & ~n4216;
  assign n4218 = ~n4198 & ~n4217;
  assign n4219 = ~n4197 & ~n4218;
  assign n4220 = ~n4196 & ~n4219;
  assign n4221 = ~n4195 & ~n4220;
  assign n4222 = ~n4194 & ~n4221;
  assign n4223 = ~pi103 & pi119;
  assign n4224 = pi103 & ~pi119;
  assign n4225 = ~pi104 & pi120;
  assign n4226 = pi104 & ~pi120;
  assign n4227 = ~pi105 & pi121;
  assign n4228 = pi105 & ~pi121;
  assign n4229 = ~pi106 & pi122;
  assign n4230 = pi106 & ~pi122;
  assign n4231 = ~pi107 & pi123;
  assign n4232 = pi107 & ~pi123;
  assign n4233 = ~pi108 & pi124;
  assign n4234 = pi108 & ~pi124;
  assign n4235 = pi110 & ~pi126;
  assign n4236 = pi109 & ~pi125;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~pi109 & pi125;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = ~n4234 & ~n4239;
  assign n4241 = ~n4233 & ~n4240;
  assign n4242 = ~n4232 & ~n4241;
  assign n4243 = ~n4231 & ~n4242;
  assign n4244 = ~n4230 & ~n4243;
  assign n4245 = ~n4229 & ~n4244;
  assign n4246 = ~n4228 & ~n4245;
  assign n4247 = ~n4227 & ~n4246;
  assign n4248 = ~n4226 & ~n4247;
  assign n4249 = ~n4225 & ~n4248;
  assign n4250 = ~n4224 & ~n4249;
  assign n4251 = ~n4223 & ~n4250;
  assign n4252 = ~n4222 & ~n4251;
  assign n4253 = n4193 & n4252;
  assign n4254 = ~pi103 & pi151;
  assign n4255 = pi105 & ~pi153;
  assign n4256 = ~pi106 & pi154;
  assign n4257 = pi106 & ~pi154;
  assign n4258 = ~pi107 & pi155;
  assign n4259 = pi107 & ~pi155;
  assign n4260 = ~pi108 & pi156;
  assign n4261 = pi108 & ~pi156;
  assign n4262 = pi110 & ~pi158;
  assign n4263 = pi109 & ~pi157;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = ~pi109 & pi157;
  assign n4266 = ~n4264 & ~n4265;
  assign n4267 = ~n4261 & ~n4266;
  assign n4268 = ~n4260 & ~n4267;
  assign n4269 = ~n4259 & ~n4268;
  assign n4270 = ~n4258 & ~n4269;
  assign n4271 = ~n4257 & ~n4270;
  assign n4272 = ~n4256 & ~n4271;
  assign n4273 = ~n4255 & ~n4272;
  assign n4274 = ~pi105 & pi153;
  assign n4275 = ~pi104 & pi152;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n4273 & n4276;
  assign n4278 = pi103 & ~pi151;
  assign n4279 = pi104 & ~pi152;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = ~n4277 & n4280;
  assign n4282 = ~n4254 & ~n4281;
  assign n4283 = ~pi103 & pi223;
  assign n4284 = pi105 & ~pi225;
  assign n4285 = ~pi106 & pi226;
  assign n4286 = pi106 & ~pi226;
  assign n4287 = ~pi107 & pi227;
  assign n4288 = pi107 & ~pi227;
  assign n4289 = ~pi108 & pi228;
  assign n4290 = pi108 & ~pi228;
  assign n4291 = pi110 & ~pi230;
  assign n4292 = pi109 & ~pi229;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = ~pi109 & pi229;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = ~n4290 & ~n4295;
  assign n4297 = ~n4289 & ~n4296;
  assign n4298 = ~n4288 & ~n4297;
  assign n4299 = ~n4287 & ~n4298;
  assign n4300 = ~n4286 & ~n4299;
  assign n4301 = ~n4285 & ~n4300;
  assign n4302 = ~n4284 & ~n4301;
  assign n4303 = ~pi105 & pi225;
  assign n4304 = ~pi104 & pi224;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = ~n4302 & n4305;
  assign n4307 = pi103 & ~pi223;
  assign n4308 = pi104 & ~pi224;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = ~n4306 & n4309;
  assign n4311 = ~n4283 & ~n4310;
  assign n4312 = ~n4282 & ~n4311;
  assign n4313 = ~pi103 & pi215;
  assign n4314 = pi105 & ~pi217;
  assign n4315 = ~pi106 & pi218;
  assign n4316 = pi106 & ~pi218;
  assign n4317 = ~pi107 & pi219;
  assign n4318 = pi107 & ~pi219;
  assign n4319 = ~pi108 & pi220;
  assign n4320 = pi108 & ~pi220;
  assign n4321 = pi110 & ~pi222;
  assign n4322 = pi109 & ~pi221;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~pi109 & pi221;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4320 & ~n4325;
  assign n4327 = ~n4319 & ~n4326;
  assign n4328 = ~n4318 & ~n4327;
  assign n4329 = ~n4317 & ~n4328;
  assign n4330 = ~n4316 & ~n4329;
  assign n4331 = ~n4315 & ~n4330;
  assign n4332 = ~n4314 & ~n4331;
  assign n4333 = ~pi105 & pi217;
  assign n4334 = ~pi104 & pi216;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = ~n4332 & n4335;
  assign n4337 = pi103 & ~pi215;
  assign n4338 = pi104 & ~pi216;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = ~n4336 & n4339;
  assign n4341 = ~n4313 & ~n4340;
  assign n4342 = ~pi103 & pi167;
  assign n4343 = pi105 & ~pi169;
  assign n4344 = ~pi106 & pi170;
  assign n4345 = pi106 & ~pi170;
  assign n4346 = ~pi107 & pi171;
  assign n4347 = pi107 & ~pi171;
  assign n4348 = ~pi108 & pi172;
  assign n4349 = pi108 & ~pi172;
  assign n4350 = pi110 & ~pi174;
  assign n4351 = pi109 & ~pi173;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = ~pi109 & pi173;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4349 & ~n4354;
  assign n4356 = ~n4348 & ~n4355;
  assign n4357 = ~n4347 & ~n4356;
  assign n4358 = ~n4346 & ~n4357;
  assign n4359 = ~n4345 & ~n4358;
  assign n4360 = ~n4344 & ~n4359;
  assign n4361 = ~n4343 & ~n4360;
  assign n4362 = ~pi105 & pi169;
  assign n4363 = ~pi104 & pi168;
  assign n4364 = ~n4362 & ~n4363;
  assign n4365 = ~n4361 & n4364;
  assign n4366 = pi103 & ~pi167;
  assign n4367 = pi104 & ~pi168;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = ~n4365 & n4368;
  assign n4370 = ~n4342 & ~n4369;
  assign n4371 = ~n4341 & ~n4370;
  assign n4372 = n4312 & n4371;
  assign n4373 = ~pi103 & pi271;
  assign n4374 = pi105 & ~pi273;
  assign n4375 = ~pi106 & pi274;
  assign n4376 = pi106 & ~pi274;
  assign n4377 = ~pi107 & pi275;
  assign n4378 = pi107 & ~pi275;
  assign n4379 = ~pi108 & pi276;
  assign n4380 = pi108 & ~pi276;
  assign n4381 = pi110 & ~pi278;
  assign n4382 = pi109 & ~pi277;
  assign n4383 = ~n4381 & ~n4382;
  assign n4384 = ~pi109 & pi277;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~n4380 & ~n4385;
  assign n4387 = ~n4379 & ~n4386;
  assign n4388 = ~n4378 & ~n4387;
  assign n4389 = ~n4377 & ~n4388;
  assign n4390 = ~n4376 & ~n4389;
  assign n4391 = ~n4375 & ~n4390;
  assign n4392 = ~n4374 & ~n4391;
  assign n4393 = ~pi105 & pi273;
  assign n4394 = ~pi104 & pi272;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4392 & n4395;
  assign n4397 = pi103 & ~pi271;
  assign n4398 = pi104 & ~pi272;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4396 & n4399;
  assign n4401 = ~n4373 & ~n4400;
  assign n4402 = ~pi103 & pi255;
  assign n4403 = pi105 & ~pi257;
  assign n4404 = ~pi106 & pi258;
  assign n4405 = pi106 & ~pi258;
  assign n4406 = ~pi107 & pi259;
  assign n4407 = pi107 & ~pi259;
  assign n4408 = ~pi108 & pi260;
  assign n4409 = pi108 & ~pi260;
  assign n4410 = pi110 & ~pi262;
  assign n4411 = pi109 & ~pi261;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = ~pi109 & pi261;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = ~n4409 & ~n4414;
  assign n4416 = ~n4408 & ~n4415;
  assign n4417 = ~n4407 & ~n4416;
  assign n4418 = ~n4406 & ~n4417;
  assign n4419 = ~n4405 & ~n4418;
  assign n4420 = ~n4404 & ~n4419;
  assign n4421 = ~n4403 & ~n4420;
  assign n4422 = ~pi105 & pi257;
  assign n4423 = ~pi104 & pi256;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~n4421 & n4424;
  assign n4426 = pi103 & ~pi255;
  assign n4427 = pi104 & ~pi256;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~n4425 & n4428;
  assign n4430 = ~n4402 & ~n4429;
  assign n4431 = ~n4401 & ~n4430;
  assign n4432 = ~pi103 & pi263;
  assign n4433 = pi105 & ~pi265;
  assign n4434 = ~pi106 & pi266;
  assign n4435 = pi106 & ~pi266;
  assign n4436 = ~pi107 & pi267;
  assign n4437 = pi107 & ~pi267;
  assign n4438 = ~pi108 & pi268;
  assign n4439 = pi108 & ~pi268;
  assign n4440 = pi110 & ~pi270;
  assign n4441 = pi109 & ~pi269;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~pi109 & pi269;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4439 & ~n4444;
  assign n4446 = ~n4438 & ~n4445;
  assign n4447 = ~n4437 & ~n4446;
  assign n4448 = ~n4436 & ~n4447;
  assign n4449 = ~n4435 & ~n4448;
  assign n4450 = ~n4434 & ~n4449;
  assign n4451 = ~n4433 & ~n4450;
  assign n4452 = ~pi105 & pi265;
  assign n4453 = ~pi104 & pi264;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~n4451 & n4454;
  assign n4456 = pi103 & ~pi263;
  assign n4457 = pi104 & ~pi264;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = ~n4455 & n4458;
  assign n4460 = ~n4432 & ~n4459;
  assign n4461 = ~pi103 & pi247;
  assign n4462 = pi105 & ~pi249;
  assign n4463 = ~pi106 & pi250;
  assign n4464 = pi106 & ~pi250;
  assign n4465 = ~pi107 & pi251;
  assign n4466 = pi107 & ~pi251;
  assign n4467 = ~pi108 & pi252;
  assign n4468 = pi108 & ~pi252;
  assign n4469 = pi110 & ~pi254;
  assign n4470 = pi109 & ~pi253;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = ~pi109 & pi253;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = ~n4468 & ~n4473;
  assign n4475 = ~n4467 & ~n4474;
  assign n4476 = ~n4466 & ~n4475;
  assign n4477 = ~n4465 & ~n4476;
  assign n4478 = ~n4464 & ~n4477;
  assign n4479 = ~n4463 & ~n4478;
  assign n4480 = ~n4462 & ~n4479;
  assign n4481 = ~pi105 & pi249;
  assign n4482 = ~pi104 & pi248;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = ~n4480 & n4483;
  assign n4485 = pi103 & ~pi247;
  assign n4486 = pi104 & ~pi248;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~n4484 & n4487;
  assign n4489 = ~n4461 & ~n4488;
  assign n4490 = ~n4460 & ~n4489;
  assign n4491 = n4431 & n4490;
  assign n4492 = n4372 & n4491;
  assign n4493 = ~pi103 & pi159;
  assign n4494 = pi103 & ~pi159;
  assign n4495 = ~pi104 & pi160;
  assign n4496 = pi104 & ~pi160;
  assign n4497 = ~pi105 & pi161;
  assign n4498 = pi105 & ~pi161;
  assign n4499 = ~pi106 & pi162;
  assign n4500 = pi106 & ~pi162;
  assign n4501 = ~pi107 & pi163;
  assign n4502 = pi107 & ~pi163;
  assign n4503 = ~pi108 & pi164;
  assign n4504 = pi108 & ~pi164;
  assign n4505 = pi110 & ~pi166;
  assign n4506 = pi109 & ~pi165;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = ~pi109 & pi165;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = ~n4504 & ~n4509;
  assign n4511 = ~n4503 & ~n4510;
  assign n4512 = ~n4502 & ~n4511;
  assign n4513 = ~n4501 & ~n4512;
  assign n4514 = ~n4500 & ~n4513;
  assign n4515 = ~n4499 & ~n4514;
  assign n4516 = ~n4498 & ~n4515;
  assign n4517 = ~n4497 & ~n4516;
  assign n4518 = ~n4496 & ~n4517;
  assign n4519 = ~n4495 & ~n4518;
  assign n4520 = ~n4494 & ~n4519;
  assign n4521 = ~n4493 & ~n4520;
  assign n4522 = ~pi103 & pi135;
  assign n4523 = pi105 & ~pi137;
  assign n4524 = ~pi106 & pi138;
  assign n4525 = pi106 & ~pi138;
  assign n4526 = ~pi107 & pi139;
  assign n4527 = pi107 & ~pi139;
  assign n4528 = ~pi108 & pi140;
  assign n4529 = pi108 & ~pi140;
  assign n4530 = pi110 & ~pi142;
  assign n4531 = pi109 & ~pi141;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~pi109 & pi141;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4529 & ~n4534;
  assign n4536 = ~n4528 & ~n4535;
  assign n4537 = ~n4527 & ~n4536;
  assign n4538 = ~n4526 & ~n4537;
  assign n4539 = ~n4525 & ~n4538;
  assign n4540 = ~n4524 & ~n4539;
  assign n4541 = ~n4523 & ~n4540;
  assign n4542 = ~pi105 & pi137;
  assign n4543 = ~pi104 & pi136;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = ~n4541 & n4544;
  assign n4546 = pi103 & ~pi135;
  assign n4547 = pi104 & ~pi136;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4545 & n4548;
  assign n4550 = ~n4522 & ~n4549;
  assign n4551 = ~pi103 & pi199;
  assign n4552 = pi105 & ~pi201;
  assign n4553 = ~pi106 & pi202;
  assign n4554 = pi106 & ~pi202;
  assign n4555 = ~pi107 & pi203;
  assign n4556 = pi107 & ~pi203;
  assign n4557 = ~pi108 & pi204;
  assign n4558 = pi108 & ~pi204;
  assign n4559 = pi110 & ~pi206;
  assign n4560 = pi109 & ~pi205;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~pi109 & pi205;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = ~n4558 & ~n4563;
  assign n4565 = ~n4557 & ~n4564;
  assign n4566 = ~n4556 & ~n4565;
  assign n4567 = ~n4555 & ~n4566;
  assign n4568 = ~n4554 & ~n4567;
  assign n4569 = ~n4553 & ~n4568;
  assign n4570 = ~n4552 & ~n4569;
  assign n4571 = ~pi105 & pi201;
  assign n4572 = ~pi104 & pi200;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = ~n4570 & n4573;
  assign n4575 = pi103 & ~pi199;
  assign n4576 = pi104 & ~pi200;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = ~n4574 & n4577;
  assign n4579 = ~n4551 & ~n4578;
  assign n4580 = ~pi103 & pi207;
  assign n4581 = pi105 & ~pi209;
  assign n4582 = ~pi106 & pi210;
  assign n4583 = pi106 & ~pi210;
  assign n4584 = ~pi107 & pi211;
  assign n4585 = pi107 & ~pi211;
  assign n4586 = ~pi108 & pi212;
  assign n4587 = pi108 & ~pi212;
  assign n4588 = pi110 & ~pi214;
  assign n4589 = pi109 & ~pi213;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = ~pi109 & pi213;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = ~n4587 & ~n4592;
  assign n4594 = ~n4586 & ~n4593;
  assign n4595 = ~n4585 & ~n4594;
  assign n4596 = ~n4584 & ~n4595;
  assign n4597 = ~n4583 & ~n4596;
  assign n4598 = ~n4582 & ~n4597;
  assign n4599 = ~n4581 & ~n4598;
  assign n4600 = ~pi105 & pi209;
  assign n4601 = ~pi104 & pi208;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4599 & n4602;
  assign n4604 = pi103 & ~pi207;
  assign n4605 = pi104 & ~pi208;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = ~n4603 & n4606;
  assign n4608 = ~n4580 & ~n4607;
  assign n4609 = ~n4579 & ~n4608;
  assign n4610 = ~n4550 & n4609;
  assign n4611 = ~n4521 & n4610;
  assign n4612 = n4492 & n4611;
  assign n4613 = pi009 & ~n501;
  assign n4614 = n2311 & n4613;
  assign n4615 = n3813 & n4614;
  assign n4616 = n3811 & n4615;
  assign n4617 = ~n2306 & n4616;
  assign n4618 = n3819 & n4617;
  assign n4619 = n3823 & n4618;
  assign n4620 = ~pi103 & pi127;
  assign n4621 = pi105 & ~pi129;
  assign n4622 = ~pi106 & pi130;
  assign n4623 = pi106 & ~pi130;
  assign n4624 = ~pi107 & pi131;
  assign n4625 = pi107 & ~pi131;
  assign n4626 = ~pi108 & pi132;
  assign n4627 = pi108 & ~pi132;
  assign n4628 = pi110 & ~pi134;
  assign n4629 = pi109 & ~pi133;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = ~pi109 & pi133;
  assign n4632 = ~n4630 & ~n4631;
  assign n4633 = ~n4627 & ~n4632;
  assign n4634 = ~n4626 & ~n4633;
  assign n4635 = ~n4625 & ~n4634;
  assign n4636 = ~n4624 & ~n4635;
  assign n4637 = ~n4623 & ~n4636;
  assign n4638 = ~n4622 & ~n4637;
  assign n4639 = ~n4621 & ~n4638;
  assign n4640 = ~pi105 & pi129;
  assign n4641 = ~pi104 & pi128;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n4639 & n4642;
  assign n4644 = pi103 & ~pi127;
  assign n4645 = pi104 & ~pi128;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4643 & n4646;
  assign n4648 = ~n4620 & ~n4647;
  assign n4649 = ~pi103 & pi183;
  assign n4650 = pi105 & ~pi185;
  assign n4651 = ~pi106 & pi186;
  assign n4652 = pi106 & ~pi186;
  assign n4653 = ~pi107 & pi187;
  assign n4654 = pi107 & ~pi187;
  assign n4655 = ~pi108 & pi188;
  assign n4656 = pi108 & ~pi188;
  assign n4657 = pi110 & ~pi190;
  assign n4658 = pi109 & ~pi189;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~pi109 & pi189;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = ~n4656 & ~n4661;
  assign n4663 = ~n4655 & ~n4662;
  assign n4664 = ~n4654 & ~n4663;
  assign n4665 = ~n4653 & ~n4664;
  assign n4666 = ~n4652 & ~n4665;
  assign n4667 = ~n4651 & ~n4666;
  assign n4668 = ~n4650 & ~n4667;
  assign n4669 = ~pi105 & pi185;
  assign n4670 = ~pi104 & pi184;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = ~n4668 & n4671;
  assign n4673 = pi103 & ~pi183;
  assign n4674 = pi104 & ~pi184;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = ~n4672 & n4675;
  assign n4677 = ~n4649 & ~n4676;
  assign n4678 = ~n4648 & ~n4677;
  assign n4679 = ~pi103 & pi239;
  assign n4680 = pi105 & ~pi241;
  assign n4681 = ~pi106 & pi242;
  assign n4682 = pi106 & ~pi242;
  assign n4683 = ~pi107 & pi243;
  assign n4684 = pi107 & ~pi243;
  assign n4685 = ~pi108 & pi244;
  assign n4686 = pi108 & ~pi244;
  assign n4687 = pi110 & ~pi246;
  assign n4688 = pi109 & ~pi245;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~pi109 & pi245;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = ~n4686 & ~n4691;
  assign n4693 = ~n4685 & ~n4692;
  assign n4694 = ~n4684 & ~n4693;
  assign n4695 = ~n4683 & ~n4694;
  assign n4696 = ~n4682 & ~n4695;
  assign n4697 = ~n4681 & ~n4696;
  assign n4698 = ~n4680 & ~n4697;
  assign n4699 = ~pi105 & pi241;
  assign n4700 = ~pi104 & pi240;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~n4698 & n4701;
  assign n4703 = pi103 & ~pi239;
  assign n4704 = pi104 & ~pi240;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = ~n4702 & n4705;
  assign n4707 = ~n4679 & ~n4706;
  assign n4708 = ~pi103 & pi231;
  assign n4709 = pi105 & ~pi233;
  assign n4710 = ~pi106 & pi234;
  assign n4711 = pi106 & ~pi234;
  assign n4712 = ~pi107 & pi235;
  assign n4713 = pi107 & ~pi235;
  assign n4714 = ~pi108 & pi236;
  assign n4715 = pi108 & ~pi236;
  assign n4716 = pi110 & ~pi238;
  assign n4717 = pi109 & ~pi237;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~pi109 & pi237;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4715 & ~n4720;
  assign n4722 = ~n4714 & ~n4721;
  assign n4723 = ~n4713 & ~n4722;
  assign n4724 = ~n4712 & ~n4723;
  assign n4725 = ~n4711 & ~n4724;
  assign n4726 = ~n4710 & ~n4725;
  assign n4727 = ~n4709 & ~n4726;
  assign n4728 = ~pi105 & pi233;
  assign n4729 = ~pi104 & pi232;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = ~n4727 & n4730;
  assign n4732 = pi103 & ~pi231;
  assign n4733 = pi104 & ~pi232;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = ~n4731 & n4734;
  assign n4736 = ~n4708 & ~n4735;
  assign n4737 = ~n4707 & ~n4736;
  assign n4738 = n4678 & n4737;
  assign n4739 = ~pi103 & pi111;
  assign n4740 = pi105 & ~pi113;
  assign n4741 = ~pi106 & pi114;
  assign n4742 = pi106 & ~pi114;
  assign n4743 = ~pi107 & pi115;
  assign n4744 = pi107 & ~pi115;
  assign n4745 = ~pi108 & pi116;
  assign n4746 = pi108 & ~pi116;
  assign n4747 = pi110 & ~pi118;
  assign n4748 = pi109 & ~pi117;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~pi109 & pi117;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4746 & ~n4751;
  assign n4753 = ~n4745 & ~n4752;
  assign n4754 = ~n4744 & ~n4753;
  assign n4755 = ~n4743 & ~n4754;
  assign n4756 = ~n4742 & ~n4755;
  assign n4757 = ~n4741 & ~n4756;
  assign n4758 = ~n4740 & ~n4757;
  assign n4759 = ~pi105 & pi113;
  assign n4760 = ~pi104 & pi112;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = ~n4758 & n4761;
  assign n4763 = pi103 & ~pi111;
  assign n4764 = pi104 & ~pi112;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = ~n4762 & n4765;
  assign n4767 = ~n4739 & ~n4766;
  assign n4768 = ~n1493 & ~n4767;
  assign n4769 = n3808 & n4768;
  assign n4770 = n4738 & n4769;
  assign n4771 = n4619 & n4770;
  assign n4772 = n4612 & n4771;
  assign n4773 = n4253 & n4772;
  assign n4774 = ~n4134 & n4773;
  assign n4775 = ~n3224 & ~n3940;
  assign n4776 = ~n1835 & ~n2242;
  assign n4777 = ~n3095 & n4776;
  assign n4778 = ~n3997 & n4777;
  assign n4779 = ~n875 & ~n1372;
  assign n4780 = ~n2243 & n4779;
  assign n4781 = ~n3104 & n4780;
  assign n4782 = ~n3971 & n4781;
  assign n4783 = ~n4778 & ~n4782;
  assign n4784 = ~n4775 & n4783;
  assign n4785 = n4774 & n4784;
  assign n4786 = ~n1432 & ~n1493;
  assign n4787 = n3808 & n4786;
  assign n4788 = ~n2691 & ~n3254;
  assign n4789 = ~n4766 & n4788;
  assign n4790 = n2219 & n3812;
  assign n4791 = pi010 & ~n501;
  assign n4792 = ~n504 & ~n969;
  assign n4793 = n4791 & n4792;
  assign n4794 = n4790 & n4793;
  assign n4795 = ~n2664 & ~n3285;
  assign n4796 = ~n3227 & ~n4739;
  assign n4797 = n4795 & n4796;
  assign n4798 = ~n1404 & ~n1435;
  assign n4799 = n3810 & n4798;
  assign n4800 = n4797 & n4799;
  assign n4801 = n4794 & n4800;
  assign n4802 = ~n996 & n4801;
  assign n4803 = ~n2306 & n4802;
  assign n4804 = n3819 & n4803;
  assign n4805 = n4789 & n4804;
  assign n4806 = n3823 & n4805;
  assign n4807 = n4787 & n4806;
  assign n4808 = ~n4785 & ~n4807;
  assign n4809 = ~n4132 & n4808;
  assign po005 = n4129 | ~n4809;
  assign n4811 = ~n3255 & ~n3940;
  assign n4812 = ~n4001 & n4811;
  assign n4813 = n3948 & n4770;
  assign n4814 = n4612 & n4813;
  assign n4815 = n4253 & n4814;
  assign n4816 = ~n4134 & n4815;
  assign n4817 = n4784 & n4816;
  assign n4818 = ~n4767 & ~n4817;
  assign n4819 = ~n2692 & ~n3066;
  assign n4820 = ~n3983 & n4819;
  assign n4821 = ~n4024 & n4820;
  assign n4822 = ~n4818 & ~n4821;
  assign n4823 = ~n4812 & n4822;
  assign n4824 = n1680 & n3086;
  assign n4825 = n3883 & n4824;
  assign n4826 = n3882 & n4825;
  assign n4827 = n1989 & n3080;
  assign n4828 = n3085 & n3088;
  assign n4829 = n1928 & n4828;
  assign n4830 = n4827 & n4829;
  assign n4831 = n4826 & n4830;
  assign n4832 = ~n4025 & n4831;
  assign n4833 = ~n2242 & n4832;
  assign n4834 = ~n3095 & n4833;
  assign n4835 = ~n3997 & n4834;
  assign n4836 = ~n4003 & n4835;
  assign n4837 = n4044 & n4836;
  assign n4838 = ~n1433 & ~n2242;
  assign n4839 = ~n3095 & n4838;
  assign n4840 = ~n3997 & n4839;
  assign n4841 = ~n4837 & n4840;
  assign n4842 = ~n4003 & ~n4069;
  assign n4843 = ~n4068 & ~n4070;
  assign n4844 = n4842 & n4843;
  assign n4845 = n3932 & ~n4844;
  assign n4846 = n3812 & n4798;
  assign n4847 = n2246 & n4792;
  assign n4848 = n4846 & n4847;
  assign n4849 = ~n2664 & ~n3227;
  assign n4850 = ~n4739 & n4849;
  assign n4851 = n3942 & n4850;
  assign n4852 = n4848 & n4851;
  assign n4853 = ~n996 & n4852;
  assign n4854 = ~n2306 & n4853;
  assign n4855 = n3819 & n4854;
  assign n4856 = n4789 & n4855;
  assign n4857 = n3823 & n4856;
  assign n4858 = n4787 & n4857;
  assign n4859 = ~n4845 & ~n4858;
  assign n4860 = ~n4841 & n4859;
  assign n4861 = n843 & n1369;
  assign n4862 = n720 & n4861;
  assign n4863 = n4048 & n4862;
  assign n4864 = ~n4047 & n4863;
  assign n4865 = n3831 & n4864;
  assign n4866 = ~n3104 & n4865;
  assign n4867 = ~n3971 & n4866;
  assign n4868 = ~n4003 & n4867;
  assign n4869 = ~n4046 & ~n4059;
  assign n4870 = ~n4058 & ~n4060;
  assign n4871 = n4869 & n4870;
  assign n4872 = n4868 & n4871;
  assign n4873 = ~n997 & ~n1372;
  assign n4874 = ~n2243 & n4873;
  assign n4875 = ~n3104 & n4874;
  assign n4876 = ~n3971 & n4875;
  assign n4877 = ~n4872 & n4876;
  assign n4878 = ~po149 & ~n4128;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = n4860 & n4879;
  assign n4881 = n4823 & n4880;
  assign n4882 = ~n4024 & n4134;
  assign n4883 = n4782 & ~n4872;
  assign n4884 = n4778 & ~n4837;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = ~n4882 & n4885;
  assign n4887 = n4767 & ~n4858;
  assign n4888 = ~n4192 & ~n4222;
  assign n4889 = ~n4251 & n4888;
  assign n4890 = n4491 & n4738;
  assign n4891 = n4372 & n4610;
  assign n4892 = ~n4163 & ~n4521;
  assign n4893 = n4891 & n4892;
  assign n4894 = n4890 & n4893;
  assign n4895 = n4889 & n4894;
  assign n4896 = ~n4887 & n4895;
  assign n4897 = ~n4817 & n4896;
  assign n4898 = ~n4845 & n4897;
  assign n4899 = ~n4001 & n4775;
  assign n4900 = ~n4878 & ~n4899;
  assign n4901 = n4898 & n4900;
  assign n4902 = n4886 & n4901;
  assign n4903 = ~n4024 & n4068;
  assign n4904 = n3932 & ~n4003;
  assign n4905 = ~n4844 & n4904;
  assign n4906 = ~n4903 & n4905;
  assign n4907 = n4070 & ~n4837;
  assign n4908 = n4069 & ~n4872;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = n4906 & n4909;
  assign n4911 = n875 & ~n4817;
  assign n4912 = n4046 & ~n4837;
  assign n4913 = ~n4024 & n4059;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = ~n4911 & n4914;
  assign n4916 = n4058 & ~n4844;
  assign n4917 = n997 & ~n4858;
  assign n4918 = n1056 & n1176;
  assign n4919 = ~n1208 & n4918;
  assign n4920 = ~n750 & ~n1238;
  assign n4921 = n4919 & n4920;
  assign n4922 = ~n1086 & ~n1328;
  assign n4923 = ~n1299 & ~n1357;
  assign n4924 = n4922 & n4923;
  assign n4925 = ~n1270 & n4924;
  assign n4926 = n4921 & n4925;
  assign n4927 = ~n657 & ~n688;
  assign n4928 = ~n718 & n4927;
  assign n4929 = ~n780 & ~n811;
  assign n4930 = ~n627 & ~n841;
  assign n4931 = n4929 & n4930;
  assign n4932 = n4928 & n4931;
  assign n4933 = n4926 & n4932;
  assign n4934 = ~n4917 & n4933;
  assign n4935 = ~n1372 & n4934;
  assign n4936 = ~n2243 & n4935;
  assign n4937 = ~n3104 & n4936;
  assign n4938 = ~n3837 & n4937;
  assign n4939 = ~n3971 & n4938;
  assign n4940 = ~n4872 & n4939;
  assign n4941 = ~n4916 & n4940;
  assign n4942 = n4047 & ~n4128;
  assign n4943 = ~n4001 & n4060;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = n4941 & n4944;
  assign n4946 = n4915 & n4945;
  assign n4947 = ~n4024 & n4038;
  assign n4948 = n4039 & ~n4872;
  assign n4949 = n1835 & ~n4817;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4947 & n4950;
  assign n4952 = n4042 & ~n4844;
  assign n4953 = n1433 & ~n4858;
  assign n4954 = n3069 & n3075;
  assign n4955 = n3068 & n3072;
  assign n4956 = n2051 & n4026;
  assign n4957 = n4955 & n4956;
  assign n4958 = n4954 & n4957;
  assign n4959 = ~n1804 & n1989;
  assign n4960 = n1928 & n2255;
  assign n4961 = n4959 & n4960;
  assign n4962 = n4958 & n4961;
  assign n4963 = ~n4953 & n4962;
  assign n4964 = ~n2242 & n4963;
  assign n4965 = ~n3095 & n4964;
  assign n4966 = ~n3997 & n4965;
  assign n4967 = ~n4003 & n4966;
  assign n4968 = ~n4837 & n4967;
  assign n4969 = ~n4952 & n4968;
  assign n4970 = n4025 & ~n4128;
  assign n4971 = ~n4001 & n4041;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = n4969 & n4972;
  assign n4974 = n4951 & n4973;
  assign n4975 = n4017 & ~n4837;
  assign n4976 = n2905 & ~n4817;
  assign n4977 = n4020 & ~n4872;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = ~n4975 & n4978;
  assign n4980 = n4021 & ~n4844;
  assign n4981 = n2692 & ~n4858;
  assign n4982 = ~n2934 & ~n3053;
  assign n4983 = ~n2876 & n4982;
  assign n4984 = ~n2722 & n3838;
  assign n4985 = n3851 & n4984;
  assign n4986 = n4009 & n4985;
  assign n4987 = n4007 & n4986;
  assign n4988 = n4983 & n4987;
  assign n4989 = ~n4981 & n4988;
  assign n4990 = ~n3066 & n4989;
  assign n4991 = ~n3983 & n4990;
  assign n4992 = ~n4003 & n4991;
  assign n4993 = ~n4024 & n4992;
  assign n4994 = ~n4980 & n4993;
  assign n4995 = n4004 & ~n4128;
  assign n4996 = ~n4001 & n4018;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = n4994 & n4997;
  assign n4999 = n4979 & n4998;
  assign n5000 = ~n4974 & ~n4999;
  assign n5001 = ~n4946 & n5000;
  assign n5002 = n2454 & n2632;
  assign n5003 = ~pi005 & ~n2363;
  assign n5004 = n2573 & n5003;
  assign n5005 = n5002 & n5004;
  assign n5006 = ~n2663 & ~n2722;
  assign n5007 = n2843 & n5006;
  assign n5008 = n2513 & n2784;
  assign n5009 = n5007 & n5008;
  assign n5010 = n4009 & n5009;
  assign n5011 = n5005 & n5010;
  assign n5012 = n4983 & n5011;
  assign n5013 = ~n4981 & n5012;
  assign n5014 = ~n3066 & n5013;
  assign n5015 = ~n3983 & n5014;
  assign n5016 = ~n4003 & n5015;
  assign n5017 = ~n4024 & n5016;
  assign n5018 = ~n4980 & n5017;
  assign n5019 = n4997 & n5018;
  assign n5020 = n4979 & n5019;
  assign n5021 = ~n5001 & ~n5020;
  assign n5022 = ~n4910 & ~n5021;
  assign n5023 = n3998 & ~n4837;
  assign n5024 = n3950 & ~n4128;
  assign n5025 = n3984 & ~n4024;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = ~n5023 & n5026;
  assign n5028 = n3255 & ~n4858;
  assign n5029 = n3166 & ~n3195;
  assign n5030 = ~n3284 & n3433;
  assign n5031 = n3956 & n5030;
  assign n5032 = n3494 & n5031;
  assign n5033 = n3953 & n5032;
  assign n5034 = n5029 & n5033;
  assign n5035 = ~n5028 & n5034;
  assign n5036 = ~n3940 & n5035;
  assign n5037 = ~n4001 & n5036;
  assign n5038 = ~n4845 & n5037;
  assign n5039 = n3224 & ~n4817;
  assign n5040 = n3972 & ~n4872;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n5038 & n5041;
  assign n5043 = n5027 & n5042;
  assign n5044 = ~pi006 & ~n3864;
  assign n5045 = ~n3931 & n5044;
  assign n5046 = ~n4003 & n5045;
  assign n5047 = ~n4844 & n5046;
  assign n5048 = ~n4903 & n5047;
  assign n5049 = n4909 & n5048;
  assign n5050 = ~n4845 & n4878;
  assign n5051 = n4119 & ~n4837;
  assign n5052 = ~n4024 & n4116;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = n4124 & ~n4872;
  assign n5055 = ~n4001 & n4125;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n5053 & n5056;
  assign n5058 = n5050 & n5057;
  assign n5059 = ~n5049 & ~n5058;
  assign n5060 = ~n5043 & n5059;
  assign n5061 = ~n5022 & n5060;
  assign n5062 = n4096 & n4102;
  assign n5063 = n4094 & n4095;
  assign n5064 = n5062 & n5063;
  assign n5065 = n4089 & n4100;
  assign n5066 = n4099 & n4103;
  assign n5067 = n5065 & n5066;
  assign n5068 = n3494 & n5067;
  assign n5069 = n5064 & n5068;
  assign n5070 = n5029 & n5069;
  assign n5071 = ~n5028 & n5070;
  assign n5072 = ~n3940 & n5071;
  assign n5073 = ~n4001 & n5072;
  assign n5074 = ~n4845 & n5073;
  assign n5075 = n5041 & n5074;
  assign n5076 = n5027 & n5075;
  assign n5077 = ~n4128 & n4130;
  assign n5078 = ~n4845 & n5077;
  assign n5079 = n5057 & n5078;
  assign n5080 = ~n5076 & ~n5079;
  assign n5081 = ~n5061 & n5080;
  assign n5082 = ~n4902 & ~n5081;
  assign n5083 = ~n4401 & ~n4736;
  assign n5084 = ~n4430 & ~n4460;
  assign n5085 = n5083 & n5084;
  assign n5086 = pi009 & ~n4648;
  assign n5087 = ~n4677 & ~n4707;
  assign n5088 = n5086 & n5087;
  assign n5089 = n5085 & n5088;
  assign n5090 = ~n4370 & ~n4579;
  assign n5091 = ~n4550 & ~n4608;
  assign n5092 = n5090 & n5091;
  assign n5093 = ~n4282 & ~n4489;
  assign n5094 = ~n4311 & ~n4341;
  assign n5095 = n5093 & n5094;
  assign n5096 = n5092 & n5095;
  assign n5097 = n4892 & n5096;
  assign n5098 = n5089 & n5097;
  assign n5099 = n4889 & n5098;
  assign n5100 = ~n4887 & n5099;
  assign n5101 = ~n4817 & n5100;
  assign n5102 = ~n4845 & n5101;
  assign n5103 = n4900 & n5102;
  assign n5104 = n4886 & n5103;
  assign n5105 = ~n5082 & ~n5104;
  assign n5106 = ~n4881 & ~n5105;
  assign n5107 = pi010 & ~n4858;
  assign n5108 = ~n4845 & n5107;
  assign n5109 = ~n4841 & n5108;
  assign n5110 = n4879 & n5109;
  assign n5111 = n4823 & n5110;
  assign n5112 = ~n4251 & ~n4817;
  assign n5113 = ~pi119 & pi143;
  assign n5114 = pi119 & ~pi143;
  assign n5115 = ~pi120 & pi144;
  assign n5116 = pi120 & ~pi144;
  assign n5117 = ~pi121 & pi145;
  assign n5118 = pi121 & ~pi145;
  assign n5119 = ~pi122 & pi146;
  assign n5120 = pi122 & ~pi146;
  assign n5121 = ~pi123 & pi147;
  assign n5122 = pi123 & ~pi147;
  assign n5123 = ~pi124 & pi148;
  assign n5124 = pi124 & ~pi148;
  assign n5125 = pi126 & ~pi150;
  assign n5126 = pi125 & ~pi149;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = ~pi125 & pi149;
  assign n5129 = ~n5127 & ~n5128;
  assign n5130 = ~n5124 & ~n5129;
  assign n5131 = ~n5123 & ~n5130;
  assign n5132 = ~n5122 & ~n5131;
  assign n5133 = ~n5121 & ~n5132;
  assign n5134 = ~n5120 & ~n5133;
  assign n5135 = ~n5119 & ~n5134;
  assign n5136 = ~n5118 & ~n5135;
  assign n5137 = ~n5117 & ~n5136;
  assign n5138 = ~n5116 & ~n5137;
  assign n5139 = ~n5115 & ~n5138;
  assign n5140 = ~n5114 & ~n5139;
  assign n5141 = ~n5113 & ~n5140;
  assign n5142 = ~pi119 & pi191;
  assign n5143 = pi119 & ~pi191;
  assign n5144 = ~pi120 & pi192;
  assign n5145 = pi120 & ~pi192;
  assign n5146 = ~pi121 & pi193;
  assign n5147 = pi121 & ~pi193;
  assign n5148 = ~pi122 & pi194;
  assign n5149 = pi122 & ~pi194;
  assign n5150 = ~pi123 & pi195;
  assign n5151 = pi123 & ~pi195;
  assign n5152 = ~pi124 & pi196;
  assign n5153 = pi124 & ~pi196;
  assign n5154 = pi126 & ~pi198;
  assign n5155 = pi125 & ~pi197;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~pi125 & pi197;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = ~n5153 & ~n5158;
  assign n5160 = ~n5152 & ~n5159;
  assign n5161 = ~n5151 & ~n5160;
  assign n5162 = ~n5150 & ~n5161;
  assign n5163 = ~n5149 & ~n5162;
  assign n5164 = ~n5148 & ~n5163;
  assign n5165 = ~n5147 & ~n5164;
  assign n5166 = ~n5146 & ~n5165;
  assign n5167 = ~n5145 & ~n5166;
  assign n5168 = ~n5144 & ~n5167;
  assign n5169 = ~n5143 & ~n5168;
  assign n5170 = ~n5142 & ~n5169;
  assign n5171 = ~pi119 & pi159;
  assign n5172 = pi119 & ~pi159;
  assign n5173 = ~pi120 & pi160;
  assign n5174 = pi120 & ~pi160;
  assign n5175 = ~pi121 & pi161;
  assign n5176 = pi121 & ~pi161;
  assign n5177 = ~pi122 & pi162;
  assign n5178 = pi122 & ~pi162;
  assign n5179 = ~pi123 & pi163;
  assign n5180 = pi123 & ~pi163;
  assign n5181 = ~pi124 & pi164;
  assign n5182 = pi124 & ~pi164;
  assign n5183 = pi126 & ~pi166;
  assign n5184 = pi125 & ~pi165;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = ~pi125 & pi165;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = ~n5182 & ~n5187;
  assign n5189 = ~n5181 & ~n5188;
  assign n5190 = ~n5180 & ~n5189;
  assign n5191 = ~n5179 & ~n5190;
  assign n5192 = ~n5178 & ~n5191;
  assign n5193 = ~n5177 & ~n5192;
  assign n5194 = ~n5176 & ~n5193;
  assign n5195 = ~n5175 & ~n5194;
  assign n5196 = ~n5174 & ~n5195;
  assign n5197 = ~n5173 & ~n5196;
  assign n5198 = ~n5172 & ~n5197;
  assign n5199 = ~n5171 & ~n5198;
  assign n5200 = ~n5170 & ~n5199;
  assign n5201 = ~n5141 & n5200;
  assign n5202 = ~pi119 & pi215;
  assign n5203 = pi121 & ~pi217;
  assign n5204 = ~pi122 & pi218;
  assign n5205 = pi122 & ~pi218;
  assign n5206 = ~pi123 & pi219;
  assign n5207 = pi123 & ~pi219;
  assign n5208 = ~pi124 & pi220;
  assign n5209 = pi124 & ~pi220;
  assign n5210 = pi126 & ~pi222;
  assign n5211 = pi125 & ~pi221;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = ~pi125 & pi221;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = ~n5209 & ~n5214;
  assign n5216 = ~n5208 & ~n5215;
  assign n5217 = ~n5207 & ~n5216;
  assign n5218 = ~n5206 & ~n5217;
  assign n5219 = ~n5205 & ~n5218;
  assign n5220 = ~n5204 & ~n5219;
  assign n5221 = ~n5203 & ~n5220;
  assign n5222 = ~pi121 & pi217;
  assign n5223 = ~pi120 & pi216;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5221 & n5224;
  assign n5226 = pi119 & ~pi215;
  assign n5227 = pi120 & ~pi216;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = ~n5225 & n5228;
  assign n5230 = ~n5202 & ~n5229;
  assign n5231 = ~pi119 & pi167;
  assign n5232 = pi121 & ~pi169;
  assign n5233 = ~pi122 & pi170;
  assign n5234 = pi122 & ~pi170;
  assign n5235 = ~pi123 & pi171;
  assign n5236 = pi123 & ~pi171;
  assign n5237 = ~pi124 & pi172;
  assign n5238 = pi124 & ~pi172;
  assign n5239 = pi126 & ~pi174;
  assign n5240 = pi125 & ~pi173;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = ~pi125 & pi173;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = ~n5238 & ~n5243;
  assign n5245 = ~n5237 & ~n5244;
  assign n5246 = ~n5236 & ~n5245;
  assign n5247 = ~n5235 & ~n5246;
  assign n5248 = ~n5234 & ~n5247;
  assign n5249 = ~n5233 & ~n5248;
  assign n5250 = ~n5232 & ~n5249;
  assign n5251 = ~pi121 & pi169;
  assign n5252 = ~pi120 & pi168;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5250 & n5253;
  assign n5255 = pi119 & ~pi167;
  assign n5256 = pi120 & ~pi168;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n5254 & n5257;
  assign n5259 = ~n5231 & ~n5258;
  assign n5260 = ~n5230 & ~n5259;
  assign n5261 = ~pi119 & pi207;
  assign n5262 = pi121 & ~pi209;
  assign n5263 = ~pi122 & pi210;
  assign n5264 = pi122 & ~pi210;
  assign n5265 = ~pi123 & pi211;
  assign n5266 = pi123 & ~pi211;
  assign n5267 = ~pi124 & pi212;
  assign n5268 = pi124 & ~pi212;
  assign n5269 = pi126 & ~pi214;
  assign n5270 = pi125 & ~pi213;
  assign n5271 = ~n5269 & ~n5270;
  assign n5272 = ~pi125 & pi213;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = ~n5268 & ~n5273;
  assign n5275 = ~n5267 & ~n5274;
  assign n5276 = ~n5266 & ~n5275;
  assign n5277 = ~n5265 & ~n5276;
  assign n5278 = ~n5264 & ~n5277;
  assign n5279 = ~n5263 & ~n5278;
  assign n5280 = ~n5262 & ~n5279;
  assign n5281 = ~pi121 & pi209;
  assign n5282 = ~pi120 & pi208;
  assign n5283 = ~n5281 & ~n5282;
  assign n5284 = ~n5280 & n5283;
  assign n5285 = pi119 & ~pi207;
  assign n5286 = pi120 & ~pi208;
  assign n5287 = ~n5285 & ~n5286;
  assign n5288 = ~n5284 & n5287;
  assign n5289 = ~n5261 & ~n5288;
  assign n5290 = ~pi119 & pi151;
  assign n5291 = pi121 & ~pi153;
  assign n5292 = ~pi122 & pi154;
  assign n5293 = pi122 & ~pi154;
  assign n5294 = ~pi123 & pi155;
  assign n5295 = pi123 & ~pi155;
  assign n5296 = ~pi124 & pi156;
  assign n5297 = pi124 & ~pi156;
  assign n5298 = pi126 & ~pi158;
  assign n5299 = pi125 & ~pi157;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = ~pi125 & pi157;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5297 & ~n5302;
  assign n5304 = ~n5296 & ~n5303;
  assign n5305 = ~n5295 & ~n5304;
  assign n5306 = ~n5294 & ~n5305;
  assign n5307 = ~n5293 & ~n5306;
  assign n5308 = ~n5292 & ~n5307;
  assign n5309 = ~n5291 & ~n5308;
  assign n5310 = ~pi121 & pi153;
  assign n5311 = ~pi120 & pi152;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = ~n5309 & n5312;
  assign n5314 = pi119 & ~pi151;
  assign n5315 = pi120 & ~pi152;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = ~n5313 & n5316;
  assign n5318 = ~n5290 & ~n5317;
  assign n5319 = ~n5289 & ~n5318;
  assign n5320 = n5260 & n5319;
  assign n5321 = ~pi119 & pi271;
  assign n5322 = pi121 & ~pi273;
  assign n5323 = ~pi122 & pi274;
  assign n5324 = pi122 & ~pi274;
  assign n5325 = ~pi123 & pi275;
  assign n5326 = pi123 & ~pi275;
  assign n5327 = ~pi124 & pi276;
  assign n5328 = pi124 & ~pi276;
  assign n5329 = pi126 & ~pi278;
  assign n5330 = pi125 & ~pi277;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = ~pi125 & pi277;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5328 & ~n5333;
  assign n5335 = ~n5327 & ~n5334;
  assign n5336 = ~n5326 & ~n5335;
  assign n5337 = ~n5325 & ~n5336;
  assign n5338 = ~n5324 & ~n5337;
  assign n5339 = ~n5323 & ~n5338;
  assign n5340 = ~n5322 & ~n5339;
  assign n5341 = ~pi121 & pi273;
  assign n5342 = ~pi120 & pi272;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = ~n5340 & n5343;
  assign n5345 = pi119 & ~pi271;
  assign n5346 = pi120 & ~pi272;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = ~n5344 & n5347;
  assign n5349 = ~n5321 & ~n5348;
  assign n5350 = ~pi119 & pi239;
  assign n5351 = pi121 & ~pi241;
  assign n5352 = ~pi122 & pi242;
  assign n5353 = pi122 & ~pi242;
  assign n5354 = ~pi123 & pi243;
  assign n5355 = pi123 & ~pi243;
  assign n5356 = ~pi124 & pi244;
  assign n5357 = pi124 & ~pi244;
  assign n5358 = pi126 & ~pi246;
  assign n5359 = pi125 & ~pi245;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = ~pi125 & pi245;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = ~n5357 & ~n5362;
  assign n5364 = ~n5356 & ~n5363;
  assign n5365 = ~n5355 & ~n5364;
  assign n5366 = ~n5354 & ~n5365;
  assign n5367 = ~n5353 & ~n5366;
  assign n5368 = ~n5352 & ~n5367;
  assign n5369 = ~n5351 & ~n5368;
  assign n5370 = ~pi121 & pi241;
  assign n5371 = ~pi120 & pi240;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = ~n5369 & n5372;
  assign n5374 = pi119 & ~pi239;
  assign n5375 = pi120 & ~pi240;
  assign n5376 = ~n5374 & ~n5375;
  assign n5377 = ~n5373 & n5376;
  assign n5378 = ~n5350 & ~n5377;
  assign n5379 = ~n5349 & ~n5378;
  assign n5380 = ~pi119 & pi231;
  assign n5381 = pi121 & ~pi233;
  assign n5382 = ~pi122 & pi234;
  assign n5383 = pi122 & ~pi234;
  assign n5384 = ~pi123 & pi235;
  assign n5385 = pi123 & ~pi235;
  assign n5386 = ~pi124 & pi236;
  assign n5387 = pi124 & ~pi236;
  assign n5388 = pi126 & ~pi238;
  assign n5389 = pi125 & ~pi237;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = ~pi125 & pi237;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = ~n5387 & ~n5392;
  assign n5394 = ~n5386 & ~n5393;
  assign n5395 = ~n5385 & ~n5394;
  assign n5396 = ~n5384 & ~n5395;
  assign n5397 = ~n5383 & ~n5396;
  assign n5398 = ~n5382 & ~n5397;
  assign n5399 = ~n5381 & ~n5398;
  assign n5400 = ~pi121 & pi233;
  assign n5401 = ~pi120 & pi232;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~n5399 & n5402;
  assign n5404 = pi119 & ~pi231;
  assign n5405 = pi120 & ~pi232;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = ~n5403 & n5406;
  assign n5408 = ~n5380 & ~n5407;
  assign n5409 = ~pi119 & pi199;
  assign n5410 = pi121 & ~pi201;
  assign n5411 = ~pi122 & pi202;
  assign n5412 = pi122 & ~pi202;
  assign n5413 = ~pi123 & pi203;
  assign n5414 = pi123 & ~pi203;
  assign n5415 = ~pi124 & pi204;
  assign n5416 = pi124 & ~pi204;
  assign n5417 = pi126 & ~pi206;
  assign n5418 = pi125 & ~pi205;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = ~pi125 & pi205;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = ~n5416 & ~n5421;
  assign n5423 = ~n5415 & ~n5422;
  assign n5424 = ~n5414 & ~n5423;
  assign n5425 = ~n5413 & ~n5424;
  assign n5426 = ~n5412 & ~n5425;
  assign n5427 = ~n5411 & ~n5426;
  assign n5428 = ~n5410 & ~n5427;
  assign n5429 = ~pi121 & pi201;
  assign n5430 = ~pi120 & pi200;
  assign n5431 = ~n5429 & ~n5430;
  assign n5432 = ~n5428 & n5431;
  assign n5433 = pi119 & ~pi199;
  assign n5434 = pi120 & ~pi200;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = ~n5432 & n5435;
  assign n5437 = ~n5409 & ~n5436;
  assign n5438 = ~n5408 & ~n5437;
  assign n5439 = n5379 & n5438;
  assign n5440 = n5320 & n5439;
  assign n5441 = ~pi119 & pi175;
  assign n5442 = pi119 & ~pi175;
  assign n5443 = ~pi120 & pi176;
  assign n5444 = pi120 & ~pi176;
  assign n5445 = ~pi121 & pi177;
  assign n5446 = pi121 & ~pi177;
  assign n5447 = ~pi122 & pi178;
  assign n5448 = pi122 & ~pi178;
  assign n5449 = ~pi123 & pi179;
  assign n5450 = pi123 & ~pi179;
  assign n5451 = ~pi124 & pi180;
  assign n5452 = pi124 & ~pi180;
  assign n5453 = pi126 & ~pi182;
  assign n5454 = pi125 & ~pi181;
  assign n5455 = ~n5453 & ~n5454;
  assign n5456 = ~pi125 & pi181;
  assign n5457 = ~n5455 & ~n5456;
  assign n5458 = ~n5452 & ~n5457;
  assign n5459 = ~n5451 & ~n5458;
  assign n5460 = ~n5450 & ~n5459;
  assign n5461 = ~n5449 & ~n5460;
  assign n5462 = ~n5448 & ~n5461;
  assign n5463 = ~n5447 & ~n5462;
  assign n5464 = ~n5446 & ~n5463;
  assign n5465 = ~n5445 & ~n5464;
  assign n5466 = ~n5444 & ~n5465;
  assign n5467 = ~n5443 & ~n5466;
  assign n5468 = ~n5442 & ~n5467;
  assign n5469 = ~n5441 & ~n5468;
  assign n5470 = ~pi119 & pi135;
  assign n5471 = pi121 & ~pi137;
  assign n5472 = ~pi122 & pi138;
  assign n5473 = pi122 & ~pi138;
  assign n5474 = ~pi123 & pi139;
  assign n5475 = pi123 & ~pi139;
  assign n5476 = ~pi124 & pi140;
  assign n5477 = pi124 & ~pi140;
  assign n5478 = pi126 & ~pi142;
  assign n5479 = pi125 & ~pi141;
  assign n5480 = ~n5478 & ~n5479;
  assign n5481 = ~pi125 & pi141;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = ~n5477 & ~n5482;
  assign n5484 = ~n5476 & ~n5483;
  assign n5485 = ~n5475 & ~n5484;
  assign n5486 = ~n5474 & ~n5485;
  assign n5487 = ~n5473 & ~n5486;
  assign n5488 = ~n5472 & ~n5487;
  assign n5489 = ~n5471 & ~n5488;
  assign n5490 = ~pi121 & pi137;
  assign n5491 = ~pi120 & pi136;
  assign n5492 = ~n5490 & ~n5491;
  assign n5493 = ~n5489 & n5492;
  assign n5494 = pi119 & ~pi135;
  assign n5495 = pi120 & ~pi136;
  assign n5496 = ~n5494 & ~n5495;
  assign n5497 = ~n5493 & n5496;
  assign n5498 = ~n5470 & ~n5497;
  assign n5499 = ~pi119 & pi183;
  assign n5500 = pi121 & ~pi185;
  assign n5501 = ~pi122 & pi186;
  assign n5502 = pi122 & ~pi186;
  assign n5503 = ~pi123 & pi187;
  assign n5504 = pi123 & ~pi187;
  assign n5505 = ~pi124 & pi188;
  assign n5506 = pi124 & ~pi188;
  assign n5507 = pi126 & ~pi190;
  assign n5508 = pi125 & ~pi189;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~pi125 & pi189;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = ~n5506 & ~n5511;
  assign n5513 = ~n5505 & ~n5512;
  assign n5514 = ~n5504 & ~n5513;
  assign n5515 = ~n5503 & ~n5514;
  assign n5516 = ~n5502 & ~n5515;
  assign n5517 = ~n5501 & ~n5516;
  assign n5518 = ~n5500 & ~n5517;
  assign n5519 = ~pi121 & pi185;
  assign n5520 = ~pi120 & pi184;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = ~n5518 & n5521;
  assign n5523 = pi119 & ~pi183;
  assign n5524 = pi120 & ~pi184;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = ~n5522 & n5525;
  assign n5527 = ~n5499 & ~n5526;
  assign n5528 = ~pi119 & pi127;
  assign n5529 = pi121 & ~pi129;
  assign n5530 = ~pi122 & pi130;
  assign n5531 = pi122 & ~pi130;
  assign n5532 = ~pi123 & pi131;
  assign n5533 = pi123 & ~pi131;
  assign n5534 = ~pi124 & pi132;
  assign n5535 = pi124 & ~pi132;
  assign n5536 = pi126 & ~pi134;
  assign n5537 = pi125 & ~pi133;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~pi125 & pi133;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = ~n5535 & ~n5540;
  assign n5542 = ~n5534 & ~n5541;
  assign n5543 = ~n5533 & ~n5542;
  assign n5544 = ~n5532 & ~n5543;
  assign n5545 = ~n5531 & ~n5544;
  assign n5546 = ~n5530 & ~n5545;
  assign n5547 = ~n5529 & ~n5546;
  assign n5548 = ~pi121 & pi129;
  assign n5549 = ~pi120 & pi128;
  assign n5550 = ~n5548 & ~n5549;
  assign n5551 = ~n5547 & n5550;
  assign n5552 = pi119 & ~pi127;
  assign n5553 = pi120 & ~pi128;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = ~n5551 & n5554;
  assign n5556 = ~n5528 & ~n5555;
  assign n5557 = ~n5527 & ~n5556;
  assign n5558 = ~n5498 & n5557;
  assign n5559 = ~n5469 & n5558;
  assign n5560 = n5440 & n5559;
  assign n5561 = pi011 & ~n501;
  assign n5562 = n4792 & n5561;
  assign n5563 = n4790 & n5562;
  assign n5564 = n4800 & n5563;
  assign n5565 = ~n996 & n5564;
  assign n5566 = ~n2306 & n5565;
  assign n5567 = n3819 & n5566;
  assign n5568 = n4789 & n5567;
  assign n5569 = n3823 & n5568;
  assign n5570 = ~pi119 & pi223;
  assign n5571 = pi121 & ~pi225;
  assign n5572 = ~pi122 & pi226;
  assign n5573 = pi122 & ~pi226;
  assign n5574 = ~pi123 & pi227;
  assign n5575 = pi123 & ~pi227;
  assign n5576 = ~pi124 & pi228;
  assign n5577 = pi124 & ~pi228;
  assign n5578 = pi126 & ~pi230;
  assign n5579 = pi125 & ~pi229;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~pi125 & pi229;
  assign n5582 = ~n5580 & ~n5581;
  assign n5583 = ~n5577 & ~n5582;
  assign n5584 = ~n5576 & ~n5583;
  assign n5585 = ~n5575 & ~n5584;
  assign n5586 = ~n5574 & ~n5585;
  assign n5587 = ~n5573 & ~n5586;
  assign n5588 = ~n5572 & ~n5587;
  assign n5589 = ~n5571 & ~n5588;
  assign n5590 = ~pi121 & pi225;
  assign n5591 = ~pi120 & pi224;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = ~n5589 & n5592;
  assign n5594 = pi119 & ~pi223;
  assign n5595 = pi120 & ~pi224;
  assign n5596 = ~n5594 & ~n5595;
  assign n5597 = ~n5593 & n5596;
  assign n5598 = ~n5570 & ~n5597;
  assign n5599 = ~pi119 & pi255;
  assign n5600 = pi121 & ~pi257;
  assign n5601 = ~pi122 & pi258;
  assign n5602 = pi122 & ~pi258;
  assign n5603 = ~pi123 & pi259;
  assign n5604 = pi123 & ~pi259;
  assign n5605 = ~pi124 & pi260;
  assign n5606 = pi124 & ~pi260;
  assign n5607 = pi126 & ~pi262;
  assign n5608 = pi125 & ~pi261;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = ~pi125 & pi261;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = ~n5606 & ~n5611;
  assign n5613 = ~n5605 & ~n5612;
  assign n5614 = ~n5604 & ~n5613;
  assign n5615 = ~n5603 & ~n5614;
  assign n5616 = ~n5602 & ~n5615;
  assign n5617 = ~n5601 & ~n5616;
  assign n5618 = ~n5600 & ~n5617;
  assign n5619 = ~pi121 & pi257;
  assign n5620 = ~pi120 & pi256;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = ~n5618 & n5621;
  assign n5623 = pi119 & ~pi255;
  assign n5624 = pi120 & ~pi256;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~n5622 & n5625;
  assign n5627 = ~n5599 & ~n5626;
  assign n5628 = ~n5598 & ~n5627;
  assign n5629 = ~pi119 & pi247;
  assign n5630 = pi121 & ~pi249;
  assign n5631 = ~pi122 & pi250;
  assign n5632 = pi122 & ~pi250;
  assign n5633 = ~pi123 & pi251;
  assign n5634 = pi123 & ~pi251;
  assign n5635 = ~pi124 & pi252;
  assign n5636 = pi124 & ~pi252;
  assign n5637 = pi126 & ~pi254;
  assign n5638 = pi125 & ~pi253;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = ~pi125 & pi253;
  assign n5641 = ~n5639 & ~n5640;
  assign n5642 = ~n5636 & ~n5641;
  assign n5643 = ~n5635 & ~n5642;
  assign n5644 = ~n5634 & ~n5643;
  assign n5645 = ~n5633 & ~n5644;
  assign n5646 = ~n5632 & ~n5645;
  assign n5647 = ~n5631 & ~n5646;
  assign n5648 = ~n5630 & ~n5647;
  assign n5649 = ~pi121 & pi249;
  assign n5650 = ~pi120 & pi248;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = ~n5648 & n5651;
  assign n5653 = pi119 & ~pi247;
  assign n5654 = pi120 & ~pi248;
  assign n5655 = ~n5653 & ~n5654;
  assign n5656 = ~n5652 & n5655;
  assign n5657 = ~n5629 & ~n5656;
  assign n5658 = ~pi119 & pi263;
  assign n5659 = pi121 & ~pi265;
  assign n5660 = ~pi122 & pi266;
  assign n5661 = pi122 & ~pi266;
  assign n5662 = ~pi123 & pi267;
  assign n5663 = pi123 & ~pi267;
  assign n5664 = ~pi124 & pi268;
  assign n5665 = pi124 & ~pi268;
  assign n5666 = pi126 & ~pi270;
  assign n5667 = pi125 & ~pi269;
  assign n5668 = ~n5666 & ~n5667;
  assign n5669 = ~pi125 & pi269;
  assign n5670 = ~n5668 & ~n5669;
  assign n5671 = ~n5665 & ~n5670;
  assign n5672 = ~n5664 & ~n5671;
  assign n5673 = ~n5663 & ~n5672;
  assign n5674 = ~n5662 & ~n5673;
  assign n5675 = ~n5661 & ~n5674;
  assign n5676 = ~n5660 & ~n5675;
  assign n5677 = ~n5659 & ~n5676;
  assign n5678 = ~pi121 & pi265;
  assign n5679 = ~pi120 & pi264;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = ~n5677 & n5680;
  assign n5682 = pi119 & ~pi263;
  assign n5683 = pi120 & ~pi264;
  assign n5684 = ~n5682 & ~n5683;
  assign n5685 = ~n5681 & n5684;
  assign n5686 = ~n5658 & ~n5685;
  assign n5687 = ~n5657 & ~n5686;
  assign n5688 = n5628 & n5687;
  assign n5689 = n4787 & n5688;
  assign n5690 = n5569 & n5689;
  assign n5691 = n5560 & n5690;
  assign n5692 = n5201 & n5691;
  assign n5693 = ~n5112 & n5692;
  assign n5694 = ~n1988 & ~n2242;
  assign n5695 = ~n3095 & n5694;
  assign n5696 = ~n3997 & n5695;
  assign n5697 = ~n4837 & n5696;
  assign n5698 = ~n1328 & ~n1372;
  assign n5699 = ~n2243 & n5698;
  assign n5700 = ~n3104 & n5699;
  assign n5701 = ~n3971 & n5700;
  assign n5702 = ~n4872 & n5701;
  assign n5703 = ~n5697 & ~n5702;
  assign n5704 = ~n3195 & ~n3940;
  assign n5705 = ~n4001 & n5704;
  assign n5706 = ~n2876 & ~n3066;
  assign n5707 = ~n3983 & n5706;
  assign n5708 = ~n4024 & n5707;
  assign n5709 = ~n5705 & ~n5708;
  assign n5710 = n5703 & n5709;
  assign n5711 = n5693 & n5710;
  assign n5712 = pi012 & ~n501;
  assign n5713 = ~n969 & ~n1145;
  assign n5714 = n2311 & n5713;
  assign n5715 = n5712 & n5714;
  assign n5716 = n2308 & n3810;
  assign n5717 = ~n1404 & ~n2052;
  assign n5718 = n3812 & n5717;
  assign n5719 = n5716 & n5718;
  assign n5720 = ~n4620 & ~n5528;
  assign n5721 = n4796 & n5720;
  assign n5722 = ~n2694 & ~n3256;
  assign n5723 = n4795 & n5722;
  assign n5724 = n5721 & n5723;
  assign n5725 = n5719 & n5724;
  assign n5726 = n5715 & n5725;
  assign n5727 = ~n1172 & n5726;
  assign n5728 = ~n996 & n5727;
  assign n5729 = ~n2306 & n5728;
  assign n5730 = n3819 & n5729;
  assign n5731 = n3821 & n5730;
  assign n5732 = ~n4647 & ~n4766;
  assign n5733 = ~n5555 & n5732;
  assign n5734 = ~n2721 & ~n3283;
  assign n5735 = n4788 & n5734;
  assign n5736 = n5733 & n5735;
  assign n5737 = n5731 & n5736;
  assign n5738 = ~n1463 & n4786;
  assign n5739 = ~n2080 & ~n2110;
  assign n5740 = n3822 & n5739;
  assign n5741 = n5738 & n5740;
  assign n5742 = n5737 & n5741;
  assign n5743 = ~n5711 & ~n5742;
  assign n5744 = ~n5111 & n5743;
  assign po006 = n5106 | ~n5744;
  assign n5746 = ~n4881 & n4981;
  assign n5747 = n4995 & ~n5058;
  assign n5748 = n4996 & ~n5043;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = ~n5746 & n5749;
  assign n5751 = ~n4910 & n4980;
  assign n5752 = n3812 & n4792;
  assign n5753 = n2246 & n5752;
  assign n5754 = ~n1145 & ~n1435;
  assign n5755 = n5717 & n5754;
  assign n5756 = n3942 & n5755;
  assign n5757 = ~n4620 & ~n4739;
  assign n5758 = ~n5528 & n5757;
  assign n5759 = n4849 & n5722;
  assign n5760 = n5758 & n5759;
  assign n5761 = n5756 & n5760;
  assign n5762 = n5753 & n5761;
  assign n5763 = ~n1172 & n5762;
  assign n5764 = ~n996 & n5763;
  assign n5765 = ~n2306 & n5764;
  assign n5766 = n3819 & n5765;
  assign n5767 = n3821 & n5766;
  assign n5768 = n5736 & n5767;
  assign n5769 = n5741 & n5768;
  assign n5770 = n2722 & ~n5769;
  assign n5771 = n4009 & n4982;
  assign n5772 = n3846 & n3852;
  assign n5773 = n4005 & n5772;
  assign n5774 = n3838 & n3850;
  assign n5775 = n3849 & n3853;
  assign n5776 = n5774 & n5775;
  assign n5777 = n5773 & n5776;
  assign n5778 = n5771 & n5777;
  assign n5779 = ~n5770 & n5778;
  assign n5780 = ~n3066 & n5779;
  assign n5781 = ~n3983 & n5780;
  assign n5782 = ~n4003 & n5781;
  assign n5783 = ~n4024 & n5782;
  assign n5784 = ~n4999 & n5783;
  assign n5785 = ~n5751 & n5784;
  assign n5786 = ~n4902 & n4976;
  assign n5787 = n1056 & n1366;
  assign n5788 = ~n1208 & n5787;
  assign n5789 = n4920 & n5788;
  assign n5790 = n4925 & n5789;
  assign n5791 = n4932 & n5790;
  assign n5792 = ~n4917 & n5791;
  assign n5793 = ~n1372 & n5792;
  assign n5794 = ~n2243 & n5793;
  assign n5795 = ~n3104 & n5794;
  assign n5796 = ~n3837 & n5795;
  assign n5797 = ~n3971 & n5796;
  assign n5798 = ~n4872 & n5797;
  assign n5799 = ~n4916 & n5798;
  assign n5800 = n4944 & n5799;
  assign n5801 = n4915 & n5800;
  assign n5802 = n4977 & ~n5801;
  assign n5803 = ~n5786 & ~n5802;
  assign n5804 = n4857 & n5689;
  assign n5805 = n5560 & n5804;
  assign n5806 = n5201 & n5805;
  assign n5807 = ~n5112 & n5806;
  assign n5808 = n5710 & n5807;
  assign n5809 = n2876 & ~n5808;
  assign n5810 = ~n1403 & n1618;
  assign n5811 = n4825 & n5810;
  assign n5812 = n4829 & n4959;
  assign n5813 = n5811 & n5812;
  assign n5814 = ~n4953 & n5813;
  assign n5815 = ~n2242 & n5814;
  assign n5816 = ~n3095 & n5815;
  assign n5817 = ~n3997 & n5816;
  assign n5818 = ~n4003 & n5817;
  assign n5819 = ~n4837 & n5818;
  assign n5820 = ~n4952 & n5819;
  assign n5821 = n4972 & n5820;
  assign n5822 = n4951 & n5821;
  assign n5823 = n4975 & ~n5822;
  assign n5824 = ~n5809 & ~n5823;
  assign n5825 = n5803 & n5824;
  assign n5826 = n5785 & n5825;
  assign n5827 = n5750 & n5826;
  assign n5828 = ~n4902 & n4949;
  assign n5829 = n4970 & ~n5058;
  assign n5830 = n4948 & ~n5801;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~n5828 & n5831;
  assign n5833 = ~n4910 & n4952;
  assign n5834 = n2081 & ~n5769;
  assign n5835 = ~n1804 & ~n1958;
  assign n5836 = n1928 & n5835;
  assign n5837 = n1680 & n2051;
  assign n5838 = n2255 & n5837;
  assign n5839 = n3883 & n5810;
  assign n5840 = n5838 & n5839;
  assign n5841 = n5836 & n5840;
  assign n5842 = ~n5834 & n5841;
  assign n5843 = ~n2242 & n5842;
  assign n5844 = ~n3095 & n5843;
  assign n5845 = ~n3997 & n5844;
  assign n5846 = ~n4003 & n5845;
  assign n5847 = ~n4837 & n5846;
  assign n5848 = ~n5822 & n5847;
  assign n5849 = ~n5833 & n5848;
  assign n5850 = n4947 & ~n4999;
  assign n5851 = n4971 & ~n5043;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n4881 & n4953;
  assign n5854 = n1988 & ~n5808;
  assign n5855 = ~n5853 & ~n5854;
  assign n5856 = n5852 & n5855;
  assign n5857 = n5849 & n5856;
  assign n5858 = n5832 & n5857;
  assign n5859 = ~n4902 & n4911;
  assign n5860 = n4942 & ~n5058;
  assign n5861 = n4912 & ~n5822;
  assign n5862 = ~n5860 & ~n5861;
  assign n5863 = ~n5859 & n5862;
  assign n5864 = ~n4910 & n4916;
  assign n5865 = n1173 & ~n5769;
  assign n5866 = pi001 & ~n1144;
  assign n5867 = ~n1115 & n5866;
  assign n5868 = n1056 & n5867;
  assign n5869 = ~n1208 & n5868;
  assign n5870 = n4920 & n5869;
  assign n5871 = ~n1086 & ~n1357;
  assign n5872 = ~n1299 & n5871;
  assign n5873 = ~n1270 & n5872;
  assign n5874 = n5870 & n5873;
  assign n5875 = n4932 & n5874;
  assign n5876 = ~n5865 & n5875;
  assign n5877 = ~n1372 & n5876;
  assign n5878 = ~n2243 & n5877;
  assign n5879 = ~n3104 & n5878;
  assign n5880 = ~n3971 & n5879;
  assign n5881 = ~n4003 & n5880;
  assign n5882 = ~n4872 & n5881;
  assign n5883 = ~n5801 & n5882;
  assign n5884 = ~n5864 & n5883;
  assign n5885 = n4913 & ~n4999;
  assign n5886 = n4943 & ~n5043;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = ~n4881 & n4917;
  assign n5889 = n1328 & ~n5808;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n5887 & n5890;
  assign n5892 = n5884 & n5891;
  assign n5893 = n5863 & n5892;
  assign n5894 = ~n5858 & ~n5893;
  assign n5895 = ~n5827 & n5894;
  assign n5896 = ~n2663 & n2843;
  assign n5897 = n5008 & n5896;
  assign n5898 = n5005 & n5897;
  assign n5899 = n5771 & n5898;
  assign n5900 = ~n5770 & n5899;
  assign n5901 = ~n3066 & n5900;
  assign n5902 = ~n3983 & n5901;
  assign n5903 = ~n4003 & n5902;
  assign n5904 = ~n4024 & n5903;
  assign n5905 = ~n4999 & n5904;
  assign n5906 = ~n5751 & n5905;
  assign n5907 = n5825 & n5906;
  assign n5908 = n5750 & n5907;
  assign n5909 = n4903 & ~n4999;
  assign n5910 = ~n4903 & ~n4907;
  assign n5911 = ~n4908 & n5910;
  assign n5912 = n4905 & ~n5911;
  assign n5913 = ~n5909 & n5912;
  assign n5914 = n4907 & ~n5822;
  assign n5915 = n4908 & ~n5801;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = n5913 & n5916;
  assign n5918 = n5040 & ~n5801;
  assign n5919 = ~n4902 & n5039;
  assign n5920 = n5023 & ~n5822;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = ~n5918 & n5921;
  assign n5923 = n4845 & ~n4910;
  assign n5924 = n3284 & ~n5769;
  assign n5925 = n3166 & n3494;
  assign n5926 = n3554 & n3800;
  assign n5927 = n3434 & n3681;
  assign n5928 = n5926 & n5927;
  assign n5929 = n5925 & n5928;
  assign n5930 = ~n5924 & n5929;
  assign n5931 = ~n3940 & n5930;
  assign n5932 = ~n4001 & n5931;
  assign n5933 = ~n5043 & n5932;
  assign n5934 = ~n5923 & n5933;
  assign n5935 = n5024 & ~n5058;
  assign n5936 = ~n4881 & n5028;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = ~n4999 & n5025;
  assign n5939 = n3195 & ~n5808;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = n5937 & n5940;
  assign n5942 = n5934 & n5941;
  assign n5943 = n5922 & n5942;
  assign n5944 = ~n5917 & ~n5943;
  assign n5945 = ~n5908 & n5944;
  assign n5946 = ~n5895 & n5945;
  assign n5947 = ~n3432 & n4100;
  assign n5948 = n5066 & n5947;
  assign n5949 = n5064 & n5948;
  assign n5950 = n5925 & n5949;
  assign n5951 = ~n5924 & n5950;
  assign n5952 = ~n3940 & n5951;
  assign n5953 = ~n4001 & n5952;
  assign n5954 = ~n5043 & n5953;
  assign n5955 = ~n5923 & n5954;
  assign n5956 = n5941 & n5955;
  assign n5957 = n5922 & n5956;
  assign n5958 = n4878 & ~n5058;
  assign n5959 = ~n5923 & n5958;
  assign n5960 = n5051 & ~n5822;
  assign n5961 = n5054 & ~n5801;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5043 & n5055;
  assign n5964 = ~n4999 & n5052;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = n5962 & n5965;
  assign n5967 = n5959 & n5966;
  assign n5968 = n4067 & ~n4844;
  assign n5969 = ~n5911 & n5968;
  assign n5970 = ~n5909 & n5969;
  assign n5971 = n5916 & n5970;
  assign n5972 = ~n5967 & ~n5971;
  assign n5973 = ~n5957 & n5972;
  assign n5974 = ~n5946 & n5973;
  assign n5975 = ~pi008 & ~po149;
  assign n5976 = ~n4128 & n5975;
  assign n5977 = ~n5058 & n5976;
  assign n5978 = ~n5923 & n5977;
  assign n5979 = n5966 & n5978;
  assign n5980 = n4883 & ~n5801;
  assign n5981 = ~n4881 & n4887;
  assign n5982 = n4884 & ~n5822;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5980 & n5983;
  assign n5985 = n4648 & ~n5769;
  assign n5986 = n4888 & n4892;
  assign n5987 = n5085 & n5087;
  assign n5988 = n5096 & n5987;
  assign n5989 = n5986 & n5988;
  assign n5990 = ~n5985 & n5989;
  assign n5991 = ~n4817 & n5990;
  assign n5992 = ~n4902 & n5991;
  assign n5993 = ~n5923 & n5992;
  assign n5994 = n4882 & ~n4999;
  assign n5995 = ~n5958 & ~n5994;
  assign n5996 = n4251 & ~n5808;
  assign n5997 = n4899 & ~n5043;
  assign n5998 = ~n5996 & ~n5997;
  assign n5999 = n5995 & n5998;
  assign n6000 = n5993 & n5999;
  assign n6001 = n5984 & n6000;
  assign n6002 = ~n5979 & ~n6001;
  assign n6003 = ~n5974 & n6002;
  assign n6004 = pi009 & ~n4677;
  assign n6005 = n4737 & n6004;
  assign n6006 = n4491 & n6005;
  assign n6007 = n4891 & n6006;
  assign n6008 = n5986 & n6007;
  assign n6009 = ~n5985 & n6008;
  assign n6010 = ~n4817 & n6009;
  assign n6011 = ~n4902 & n6010;
  assign n6012 = ~n5923 & n6011;
  assign n6013 = n5999 & n6012;
  assign n6014 = n5984 & n6013;
  assign n6015 = n4877 & ~n5801;
  assign n6016 = n4818 & ~n4902;
  assign n6017 = ~n6015 & ~n6016;
  assign n6018 = n4812 & ~n5043;
  assign n6019 = n4841 & ~n5822;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n6017 & n6020;
  assign n6022 = ~n4858 & ~n4881;
  assign n6023 = ~n5923 & n6022;
  assign n6024 = n4821 & ~n4999;
  assign n6025 = ~n5958 & ~n6024;
  assign n6026 = n6023 & n6025;
  assign n6027 = n6021 & n6026;
  assign n6028 = ~n6014 & ~n6027;
  assign n6029 = ~n6003 & n6028;
  assign n6030 = n5702 & ~n5801;
  assign n6031 = ~n4999 & n5708;
  assign n6032 = n5697 & ~n5822;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = ~n6030 & n6033;
  assign n6035 = n5556 & ~n5769;
  assign n6036 = ~n5170 & ~n5469;
  assign n6037 = ~n5141 & ~n5199;
  assign n6038 = n6036 & n6037;
  assign n6039 = n5379 & n5687;
  assign n6040 = n5628 & n6039;
  assign n6041 = ~n5498 & ~n5527;
  assign n6042 = n5319 & n6041;
  assign n6043 = n5260 & n5438;
  assign n6044 = n6042 & n6043;
  assign n6045 = n6040 & n6044;
  assign n6046 = n6038 & n6045;
  assign n6047 = ~n6035 & n6046;
  assign n6048 = ~n5808 & n6047;
  assign n6049 = ~n5923 & n6048;
  assign n6050 = ~n5958 & ~n6022;
  assign n6051 = ~n5043 & n5705;
  assign n6052 = ~n4902 & n5112;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = n6050 & n6053;
  assign n6055 = n6049 & n6054;
  assign n6056 = n6034 & n6055;
  assign n6057 = ~pi010 & ~n4858;
  assign n6058 = ~n4881 & n6057;
  assign n6059 = ~n5923 & n6058;
  assign n6060 = n6025 & n6059;
  assign n6061 = n6021 & n6060;
  assign n6062 = ~n6056 & ~n6061;
  assign n6063 = ~n6029 & n6062;
  assign n6064 = ~n5349 & ~n5686;
  assign n6065 = ~n5378 & ~n5408;
  assign n6066 = n6064 & n6065;
  assign n6067 = pi011 & ~n5598;
  assign n6068 = ~n5627 & ~n5657;
  assign n6069 = n6067 & n6068;
  assign n6070 = n6066 & n6069;
  assign n6071 = ~n5318 & ~n5527;
  assign n6072 = ~n5498 & n6071;
  assign n6073 = ~n5230 & ~n5437;
  assign n6074 = ~n5259 & ~n5289;
  assign n6075 = n6073 & n6074;
  assign n6076 = n6072 & n6075;
  assign n6077 = n6070 & n6076;
  assign n6078 = n6038 & n6077;
  assign n6079 = ~n6035 & n6078;
  assign n6080 = ~n5808 & n6079;
  assign n6081 = ~n5923 & n6080;
  assign n6082 = n6054 & n6081;
  assign n6083 = n6034 & n6082;
  assign n6084 = ~n6063 & ~n6083;
  assign n6085 = ~n1173 & ~n1372;
  assign n6086 = ~n2243 & n6085;
  assign n6087 = ~n3104 & n6086;
  assign n6088 = ~n3971 & n6087;
  assign n6089 = ~n4872 & n6088;
  assign n6090 = ~n5801 & n6089;
  assign n6091 = ~n4648 & ~n4817;
  assign n6092 = ~n4902 & n6091;
  assign n6093 = ~n5556 & ~n5808;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = ~n6090 & n6094;
  assign n6096 = ~n5769 & ~n5923;
  assign n6097 = ~n5958 & n6096;
  assign n6098 = ~n2722 & ~n3066;
  assign n6099 = ~n3983 & n6098;
  assign n6100 = ~n4024 & n6099;
  assign n6101 = ~n4999 & n6100;
  assign n6102 = ~n6022 & ~n6101;
  assign n6103 = ~n2081 & ~n2242;
  assign n6104 = ~n3095 & n6103;
  assign n6105 = ~n3997 & n6104;
  assign n6106 = ~n4837 & n6105;
  assign n6107 = ~n5822 & n6106;
  assign n6108 = ~n3284 & ~n3940;
  assign n6109 = ~n4001 & n6108;
  assign n6110 = ~n5043 & n6109;
  assign n6111 = ~n6107 & ~n6110;
  assign n6112 = n6102 & n6111;
  assign n6113 = n6097 & n6112;
  assign n6114 = n6095 & n6113;
  assign n6115 = ~n6084 & ~n6114;
  assign n6116 = pi012 & ~n5769;
  assign n6117 = ~n5923 & n6116;
  assign n6118 = ~n5958 & n6117;
  assign n6119 = n6112 & n6118;
  assign n6120 = n6095 & n6119;
  assign n6121 = ~n1927 & ~n2242;
  assign n6122 = ~n3095 & n6121;
  assign n6123 = ~n3997 & n6122;
  assign n6124 = ~n4837 & n6123;
  assign n6125 = ~n5822 & n6124;
  assign n6126 = ~n1357 & ~n1372;
  assign n6127 = ~n2243 & n6126;
  assign n6128 = ~n3104 & n6127;
  assign n6129 = ~n3971 & n6128;
  assign n6130 = ~n4872 & n6129;
  assign n6131 = ~n5801 & n6130;
  assign n6132 = ~n5141 & ~n5808;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = ~n6125 & n6133;
  assign n6135 = ~n3493 & ~n3940;
  assign n6136 = ~n4001 & n6135;
  assign n6137 = ~n5043 & n6136;
  assign n6138 = n2311 & n5717;
  assign n6139 = pi014 & ~n501;
  assign n6140 = n5713 & n6139;
  assign n6141 = n6138 & n6140;
  assign n6142 = n3810 & n5722;
  assign n6143 = n3813 & n6142;
  assign n6144 = ~pi135 & pi143;
  assign n6145 = n5720 & ~n6144;
  assign n6146 = n4797 & n6145;
  assign n6147 = n6143 & n6146;
  assign n6148 = n6141 & n6147;
  assign n6149 = ~n1172 & n6148;
  assign n6150 = ~n996 & n6149;
  assign n6151 = ~n2306 & n6150;
  assign n6152 = n3819 & n6151;
  assign n6153 = n3821 & n6152;
  assign n6154 = pi137 & ~pi145;
  assign n6155 = ~pi138 & pi146;
  assign n6156 = pi138 & ~pi146;
  assign n6157 = ~pi139 & pi147;
  assign n6158 = pi139 & ~pi147;
  assign n6159 = ~pi140 & pi148;
  assign n6160 = pi140 & ~pi148;
  assign n6161 = pi142 & ~pi150;
  assign n6162 = pi141 & ~pi149;
  assign n6163 = ~n6161 & ~n6162;
  assign n6164 = ~pi141 & pi149;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = ~n6160 & ~n6165;
  assign n6167 = ~n6159 & ~n6166;
  assign n6168 = ~n6158 & ~n6167;
  assign n6169 = ~n6157 & ~n6168;
  assign n6170 = ~n6156 & ~n6169;
  assign n6171 = ~n6155 & ~n6170;
  assign n6172 = ~n6154 & ~n6171;
  assign n6173 = ~pi137 & pi145;
  assign n6174 = ~pi136 & pi144;
  assign n6175 = ~n6173 & ~n6174;
  assign n6176 = ~n6172 & n6175;
  assign n6177 = pi135 & ~pi143;
  assign n6178 = pi136 & ~pi144;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = ~n6176 & n6179;
  assign n6181 = ~n5555 & ~n6180;
  assign n6182 = n5732 & n6181;
  assign n6183 = n5735 & n6182;
  assign n6184 = n6153 & n6183;
  assign n6185 = n5741 & n6184;
  assign n6186 = ~n6137 & n6185;
  assign n6187 = ~n4222 & ~n4817;
  assign n6188 = ~n4902 & n6187;
  assign n6189 = ~n2965 & ~n3066;
  assign n6190 = ~n3983 & n6189;
  assign n6191 = ~n4024 & n6190;
  assign n6192 = ~n4999 & n6191;
  assign n6193 = ~n6188 & ~n6192;
  assign n6194 = n6186 & n6193;
  assign n6195 = n6134 & n6194;
  assign n6196 = ~pi135 & pi191;
  assign n6197 = pi135 & ~pi191;
  assign n6198 = ~pi136 & pi192;
  assign n6199 = pi136 & ~pi192;
  assign n6200 = ~pi137 & pi193;
  assign n6201 = pi137 & ~pi193;
  assign n6202 = ~pi138 & pi194;
  assign n6203 = pi138 & ~pi194;
  assign n6204 = ~pi139 & pi195;
  assign n6205 = pi139 & ~pi195;
  assign n6206 = ~pi140 & pi196;
  assign n6207 = pi140 & ~pi196;
  assign n6208 = pi142 & ~pi198;
  assign n6209 = pi141 & ~pi197;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = ~pi141 & pi197;
  assign n6212 = ~n6210 & ~n6211;
  assign n6213 = ~n6207 & ~n6212;
  assign n6214 = ~n6206 & ~n6213;
  assign n6215 = ~n6205 & ~n6214;
  assign n6216 = ~n6204 & ~n6215;
  assign n6217 = ~n6203 & ~n6216;
  assign n6218 = ~n6202 & ~n6217;
  assign n6219 = ~n6201 & ~n6218;
  assign n6220 = ~n6200 & ~n6219;
  assign n6221 = ~n6199 & ~n6220;
  assign n6222 = ~n6198 & ~n6221;
  assign n6223 = ~n6197 & ~n6222;
  assign n6224 = ~n6196 & ~n6223;
  assign n6225 = ~pi135 & pi159;
  assign n6226 = pi135 & ~pi159;
  assign n6227 = ~pi136 & pi160;
  assign n6228 = pi136 & ~pi160;
  assign n6229 = ~pi137 & pi161;
  assign n6230 = pi137 & ~pi161;
  assign n6231 = ~pi138 & pi162;
  assign n6232 = pi138 & ~pi162;
  assign n6233 = ~pi139 & pi163;
  assign n6234 = pi139 & ~pi163;
  assign n6235 = ~pi140 & pi164;
  assign n6236 = pi140 & ~pi164;
  assign n6237 = pi142 & ~pi166;
  assign n6238 = pi141 & ~pi165;
  assign n6239 = ~n6237 & ~n6238;
  assign n6240 = ~pi141 & pi165;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~n6236 & ~n6241;
  assign n6243 = ~n6235 & ~n6242;
  assign n6244 = ~n6234 & ~n6243;
  assign n6245 = ~n6233 & ~n6244;
  assign n6246 = ~n6232 & ~n6245;
  assign n6247 = ~n6231 & ~n6246;
  assign n6248 = ~n6230 & ~n6247;
  assign n6249 = ~n6229 & ~n6248;
  assign n6250 = ~n6228 & ~n6249;
  assign n6251 = ~n6227 & ~n6250;
  assign n6252 = ~n6226 & ~n6251;
  assign n6253 = ~n6225 & ~n6252;
  assign n6254 = ~pi135 & pi175;
  assign n6255 = pi135 & ~pi175;
  assign n6256 = ~pi136 & pi176;
  assign n6257 = pi136 & ~pi176;
  assign n6258 = ~pi137 & pi177;
  assign n6259 = pi137 & ~pi177;
  assign n6260 = ~pi138 & pi178;
  assign n6261 = pi138 & ~pi178;
  assign n6262 = ~pi139 & pi179;
  assign n6263 = pi139 & ~pi179;
  assign n6264 = ~pi140 & pi180;
  assign n6265 = pi140 & ~pi180;
  assign n6266 = pi142 & ~pi182;
  assign n6267 = pi141 & ~pi181;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~pi141 & pi181;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = ~n6265 & ~n6270;
  assign n6272 = ~n6264 & ~n6271;
  assign n6273 = ~n6263 & ~n6272;
  assign n6274 = ~n6262 & ~n6273;
  assign n6275 = ~n6261 & ~n6274;
  assign n6276 = ~n6260 & ~n6275;
  assign n6277 = ~n6259 & ~n6276;
  assign n6278 = ~n6258 & ~n6277;
  assign n6279 = ~n6257 & ~n6278;
  assign n6280 = ~n6256 & ~n6279;
  assign n6281 = ~n6255 & ~n6280;
  assign n6282 = ~n6254 & ~n6281;
  assign n6283 = ~n6253 & ~n6282;
  assign n6284 = ~n6224 & n6283;
  assign n6285 = ~pi135 & pi263;
  assign n6286 = pi137 & ~pi265;
  assign n6287 = ~pi138 & pi266;
  assign n6288 = pi138 & ~pi266;
  assign n6289 = ~pi139 & pi267;
  assign n6290 = pi139 & ~pi267;
  assign n6291 = ~pi140 & pi268;
  assign n6292 = pi140 & ~pi268;
  assign n6293 = pi142 & ~pi270;
  assign n6294 = pi141 & ~pi269;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = ~pi141 & pi269;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = ~n6292 & ~n6297;
  assign n6299 = ~n6291 & ~n6298;
  assign n6300 = ~n6290 & ~n6299;
  assign n6301 = ~n6289 & ~n6300;
  assign n6302 = ~n6288 & ~n6301;
  assign n6303 = ~n6287 & ~n6302;
  assign n6304 = ~n6286 & ~n6303;
  assign n6305 = ~pi137 & pi265;
  assign n6306 = ~pi136 & pi264;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = ~n6304 & n6307;
  assign n6309 = pi135 & ~pi263;
  assign n6310 = pi136 & ~pi264;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n6308 & n6311;
  assign n6313 = ~n6285 & ~n6312;
  assign n6314 = ~pi135 & pi207;
  assign n6315 = pi137 & ~pi209;
  assign n6316 = ~pi138 & pi210;
  assign n6317 = pi138 & ~pi210;
  assign n6318 = ~pi139 & pi211;
  assign n6319 = pi139 & ~pi211;
  assign n6320 = ~pi140 & pi212;
  assign n6321 = pi140 & ~pi212;
  assign n6322 = pi142 & ~pi214;
  assign n6323 = pi141 & ~pi213;
  assign n6324 = ~n6322 & ~n6323;
  assign n6325 = ~pi141 & pi213;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = ~n6321 & ~n6326;
  assign n6328 = ~n6320 & ~n6327;
  assign n6329 = ~n6319 & ~n6328;
  assign n6330 = ~n6318 & ~n6329;
  assign n6331 = ~n6317 & ~n6330;
  assign n6332 = ~n6316 & ~n6331;
  assign n6333 = ~n6315 & ~n6332;
  assign n6334 = ~pi137 & pi209;
  assign n6335 = ~pi136 & pi208;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n6333 & n6336;
  assign n6338 = pi135 & ~pi207;
  assign n6339 = pi136 & ~pi208;
  assign n6340 = ~n6338 & ~n6339;
  assign n6341 = ~n6337 & n6340;
  assign n6342 = ~n6314 & ~n6341;
  assign n6343 = ~n6313 & ~n6342;
  assign n6344 = ~pi135 & pi199;
  assign n6345 = pi137 & ~pi201;
  assign n6346 = ~pi138 & pi202;
  assign n6347 = pi138 & ~pi202;
  assign n6348 = ~pi139 & pi203;
  assign n6349 = pi139 & ~pi203;
  assign n6350 = ~pi140 & pi204;
  assign n6351 = pi140 & ~pi204;
  assign n6352 = pi142 & ~pi206;
  assign n6353 = pi141 & ~pi205;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = ~pi141 & pi205;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n6351 & ~n6356;
  assign n6358 = ~n6350 & ~n6357;
  assign n6359 = ~n6349 & ~n6358;
  assign n6360 = ~n6348 & ~n6359;
  assign n6361 = ~n6347 & ~n6360;
  assign n6362 = ~n6346 & ~n6361;
  assign n6363 = ~n6345 & ~n6362;
  assign n6364 = ~pi137 & pi201;
  assign n6365 = ~pi136 & pi200;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n6363 & n6366;
  assign n6368 = pi135 & ~pi199;
  assign n6369 = pi136 & ~pi200;
  assign n6370 = ~n6368 & ~n6369;
  assign n6371 = ~n6367 & n6370;
  assign n6372 = ~n6344 & ~n6371;
  assign n6373 = ~pi135 & pi271;
  assign n6374 = pi137 & ~pi273;
  assign n6375 = ~pi138 & pi274;
  assign n6376 = pi138 & ~pi274;
  assign n6377 = ~pi139 & pi275;
  assign n6378 = pi139 & ~pi275;
  assign n6379 = ~pi140 & pi276;
  assign n6380 = pi140 & ~pi276;
  assign n6381 = pi142 & ~pi278;
  assign n6382 = pi141 & ~pi277;
  assign n6383 = ~n6381 & ~n6382;
  assign n6384 = ~pi141 & pi277;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6380 & ~n6385;
  assign n6387 = ~n6379 & ~n6386;
  assign n6388 = ~n6378 & ~n6387;
  assign n6389 = ~n6377 & ~n6388;
  assign n6390 = ~n6376 & ~n6389;
  assign n6391 = ~n6375 & ~n6390;
  assign n6392 = ~n6374 & ~n6391;
  assign n6393 = ~pi137 & pi273;
  assign n6394 = ~pi136 & pi272;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n6392 & n6395;
  assign n6397 = pi135 & ~pi271;
  assign n6398 = pi136 & ~pi272;
  assign n6399 = ~n6397 & ~n6398;
  assign n6400 = ~n6396 & n6399;
  assign n6401 = ~n6373 & ~n6400;
  assign n6402 = ~n6372 & ~n6401;
  assign n6403 = n6343 & n6402;
  assign n6404 = ~pi135 & pi167;
  assign n6405 = pi137 & ~pi169;
  assign n6406 = ~pi138 & pi170;
  assign n6407 = pi138 & ~pi170;
  assign n6408 = ~pi139 & pi171;
  assign n6409 = pi139 & ~pi171;
  assign n6410 = ~pi140 & pi172;
  assign n6411 = pi140 & ~pi172;
  assign n6412 = pi142 & ~pi174;
  assign n6413 = pi141 & ~pi173;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = ~pi141 & pi173;
  assign n6416 = ~n6414 & ~n6415;
  assign n6417 = ~n6411 & ~n6416;
  assign n6418 = ~n6410 & ~n6417;
  assign n6419 = ~n6409 & ~n6418;
  assign n6420 = ~n6408 & ~n6419;
  assign n6421 = ~n6407 & ~n6420;
  assign n6422 = ~n6406 & ~n6421;
  assign n6423 = ~n6405 & ~n6422;
  assign n6424 = ~pi137 & pi169;
  assign n6425 = ~pi136 & pi168;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = ~n6423 & n6426;
  assign n6428 = pi135 & ~pi167;
  assign n6429 = pi136 & ~pi168;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6427 & n6430;
  assign n6432 = ~n6404 & ~n6431;
  assign n6433 = ~pi135 & pi183;
  assign n6434 = pi137 & ~pi185;
  assign n6435 = ~pi138 & pi186;
  assign n6436 = pi138 & ~pi186;
  assign n6437 = ~pi139 & pi187;
  assign n6438 = pi139 & ~pi187;
  assign n6439 = ~pi140 & pi188;
  assign n6440 = pi140 & ~pi188;
  assign n6441 = pi142 & ~pi190;
  assign n6442 = pi141 & ~pi189;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = ~pi141 & pi189;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = ~n6440 & ~n6445;
  assign n6447 = ~n6439 & ~n6446;
  assign n6448 = ~n6438 & ~n6447;
  assign n6449 = ~n6437 & ~n6448;
  assign n6450 = ~n6436 & ~n6449;
  assign n6451 = ~n6435 & ~n6450;
  assign n6452 = ~n6434 & ~n6451;
  assign n6453 = ~pi137 & pi185;
  assign n6454 = ~pi136 & pi184;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = ~n6452 & n6455;
  assign n6457 = pi135 & ~pi183;
  assign n6458 = pi136 & ~pi184;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n6456 & n6459;
  assign n6461 = ~n6433 & ~n6460;
  assign n6462 = ~n6432 & ~n6461;
  assign n6463 = n4786 & n6462;
  assign n6464 = n6403 & n6463;
  assign n6465 = ~pi135 & pi223;
  assign n6466 = pi137 & ~pi225;
  assign n6467 = ~pi138 & pi226;
  assign n6468 = pi138 & ~pi226;
  assign n6469 = ~pi139 & pi227;
  assign n6470 = pi139 & ~pi227;
  assign n6471 = ~pi140 & pi228;
  assign n6472 = pi140 & ~pi228;
  assign n6473 = pi142 & ~pi230;
  assign n6474 = pi141 & ~pi229;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~pi141 & pi229;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = ~n6472 & ~n6477;
  assign n6479 = ~n6471 & ~n6478;
  assign n6480 = ~n6470 & ~n6479;
  assign n6481 = ~n6469 & ~n6480;
  assign n6482 = ~n6468 & ~n6481;
  assign n6483 = ~n6467 & ~n6482;
  assign n6484 = ~n6466 & ~n6483;
  assign n6485 = ~pi137 & pi225;
  assign n6486 = ~pi136 & pi224;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = ~n6484 & n6487;
  assign n6489 = pi135 & ~pi223;
  assign n6490 = pi136 & ~pi224;
  assign n6491 = ~n6489 & ~n6490;
  assign n6492 = ~n6488 & n6491;
  assign n6493 = ~n6465 & ~n6492;
  assign n6494 = ~pi135 & pi239;
  assign n6495 = pi137 & ~pi241;
  assign n6496 = ~pi138 & pi242;
  assign n6497 = pi138 & ~pi242;
  assign n6498 = ~pi139 & pi243;
  assign n6499 = pi139 & ~pi243;
  assign n6500 = ~pi140 & pi244;
  assign n6501 = pi140 & ~pi244;
  assign n6502 = pi142 & ~pi246;
  assign n6503 = pi141 & ~pi245;
  assign n6504 = ~n6502 & ~n6503;
  assign n6505 = ~pi141 & pi245;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n6501 & ~n6506;
  assign n6508 = ~n6500 & ~n6507;
  assign n6509 = ~n6499 & ~n6508;
  assign n6510 = ~n6498 & ~n6509;
  assign n6511 = ~n6497 & ~n6510;
  assign n6512 = ~n6496 & ~n6511;
  assign n6513 = ~n6495 & ~n6512;
  assign n6514 = ~pi137 & pi241;
  assign n6515 = ~pi136 & pi240;
  assign n6516 = ~n6514 & ~n6515;
  assign n6517 = ~n6513 & n6516;
  assign n6518 = pi135 & ~pi239;
  assign n6519 = pi136 & ~pi240;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = ~n6517 & n6520;
  assign n6522 = ~n6494 & ~n6521;
  assign n6523 = ~n6493 & ~n6522;
  assign n6524 = ~pi135 & pi151;
  assign n6525 = pi137 & ~pi153;
  assign n6526 = ~pi138 & pi154;
  assign n6527 = pi138 & ~pi154;
  assign n6528 = ~pi139 & pi155;
  assign n6529 = pi139 & ~pi155;
  assign n6530 = ~pi140 & pi156;
  assign n6531 = pi140 & ~pi156;
  assign n6532 = pi142 & ~pi158;
  assign n6533 = pi141 & ~pi157;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = ~pi141 & pi157;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~n6531 & ~n6536;
  assign n6538 = ~n6530 & ~n6537;
  assign n6539 = ~n6529 & ~n6538;
  assign n6540 = ~n6528 & ~n6539;
  assign n6541 = ~n6527 & ~n6540;
  assign n6542 = ~n6526 & ~n6541;
  assign n6543 = ~n6525 & ~n6542;
  assign n6544 = ~pi137 & pi153;
  assign n6545 = ~pi136 & pi152;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = ~n6543 & n6546;
  assign n6548 = pi135 & ~pi151;
  assign n6549 = pi136 & ~pi152;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = ~n6547 & n6550;
  assign n6552 = ~n6524 & ~n6551;
  assign n6553 = ~n6144 & ~n6180;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n6523 & n6554;
  assign n6556 = ~pi135 & pi247;
  assign n6557 = pi137 & ~pi249;
  assign n6558 = ~pi138 & pi250;
  assign n6559 = pi138 & ~pi250;
  assign n6560 = ~pi139 & pi251;
  assign n6561 = pi139 & ~pi251;
  assign n6562 = ~pi140 & pi252;
  assign n6563 = pi140 & ~pi252;
  assign n6564 = pi142 & ~pi254;
  assign n6565 = pi141 & ~pi253;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = ~pi141 & pi253;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n6563 & ~n6568;
  assign n6570 = ~n6562 & ~n6569;
  assign n6571 = ~n6561 & ~n6570;
  assign n6572 = ~n6560 & ~n6571;
  assign n6573 = ~n6559 & ~n6572;
  assign n6574 = ~n6558 & ~n6573;
  assign n6575 = ~n6557 & ~n6574;
  assign n6576 = ~pi137 & pi249;
  assign n6577 = ~pi136 & pi248;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = ~n6575 & n6578;
  assign n6580 = pi135 & ~pi247;
  assign n6581 = pi136 & ~pi248;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n6579 & n6582;
  assign n6584 = ~n6556 & ~n6583;
  assign n6585 = ~pi135 & pi231;
  assign n6586 = pi137 & ~pi233;
  assign n6587 = ~pi138 & pi234;
  assign n6588 = pi138 & ~pi234;
  assign n6589 = ~pi139 & pi235;
  assign n6590 = pi139 & ~pi235;
  assign n6591 = ~pi140 & pi236;
  assign n6592 = pi140 & ~pi236;
  assign n6593 = pi142 & ~pi238;
  assign n6594 = pi141 & ~pi237;
  assign n6595 = ~n6593 & ~n6594;
  assign n6596 = ~pi141 & pi237;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~n6592 & ~n6597;
  assign n6599 = ~n6591 & ~n6598;
  assign n6600 = ~n6590 & ~n6599;
  assign n6601 = ~n6589 & ~n6600;
  assign n6602 = ~n6588 & ~n6601;
  assign n6603 = ~n6587 & ~n6602;
  assign n6604 = ~n6586 & ~n6603;
  assign n6605 = ~pi137 & pi233;
  assign n6606 = ~pi136 & pi232;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = ~n6604 & n6607;
  assign n6609 = pi135 & ~pi231;
  assign n6610 = pi136 & ~pi232;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = ~n6608 & n6611;
  assign n6613 = ~n6585 & ~n6612;
  assign n6614 = ~n6584 & ~n6613;
  assign n6615 = ~pi135 & pi255;
  assign n6616 = pi137 & ~pi257;
  assign n6617 = ~pi138 & pi258;
  assign n6618 = pi138 & ~pi258;
  assign n6619 = ~pi139 & pi259;
  assign n6620 = pi139 & ~pi259;
  assign n6621 = ~pi140 & pi260;
  assign n6622 = pi140 & ~pi260;
  assign n6623 = pi142 & ~pi262;
  assign n6624 = pi141 & ~pi261;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = ~pi141 & pi261;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = ~n6622 & ~n6627;
  assign n6629 = ~n6621 & ~n6628;
  assign n6630 = ~n6620 & ~n6629;
  assign n6631 = ~n6619 & ~n6630;
  assign n6632 = ~n6618 & ~n6631;
  assign n6633 = ~n6617 & ~n6632;
  assign n6634 = ~n6616 & ~n6633;
  assign n6635 = ~pi137 & pi257;
  assign n6636 = ~pi136 & pi256;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = ~n6634 & n6637;
  assign n6639 = pi135 & ~pi255;
  assign n6640 = pi136 & ~pi256;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~n6638 & n6641;
  assign n6643 = ~n6615 & ~n6642;
  assign n6644 = ~pi135 & pi215;
  assign n6645 = pi137 & ~pi217;
  assign n6646 = ~pi138 & pi218;
  assign n6647 = pi138 & ~pi218;
  assign n6648 = ~pi139 & pi219;
  assign n6649 = pi139 & ~pi219;
  assign n6650 = ~pi140 & pi220;
  assign n6651 = pi140 & ~pi220;
  assign n6652 = pi142 & ~pi222;
  assign n6653 = pi141 & ~pi221;
  assign n6654 = ~n6652 & ~n6653;
  assign n6655 = ~pi141 & pi221;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = ~n6651 & ~n6656;
  assign n6658 = ~n6650 & ~n6657;
  assign n6659 = ~n6649 & ~n6658;
  assign n6660 = ~n6648 & ~n6659;
  assign n6661 = ~n6647 & ~n6660;
  assign n6662 = ~n6646 & ~n6661;
  assign n6663 = ~n6645 & ~n6662;
  assign n6664 = ~pi137 & pi217;
  assign n6665 = ~pi136 & pi216;
  assign n6666 = ~n6664 & ~n6665;
  assign n6667 = ~n6663 & n6666;
  assign n6668 = pi135 & ~pi215;
  assign n6669 = pi136 & ~pi216;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = ~n6667 & n6670;
  assign n6672 = ~n6644 & ~n6671;
  assign n6673 = ~n6643 & ~n6672;
  assign n6674 = n6614 & n6673;
  assign n6675 = n6555 & n6674;
  assign n6676 = n6464 & n6675;
  assign n6677 = n3819 & n5734;
  assign n6678 = ~n4522 & ~n5470;
  assign n6679 = n5720 & n6678;
  assign n6680 = ~n3285 & ~n3525;
  assign n6681 = n4796 & n6680;
  assign n6682 = n6142 & n6681;
  assign n6683 = n6679 & n6682;
  assign n6684 = ~n2021 & ~n2052;
  assign n6685 = n4792 & n6684;
  assign n6686 = pi013 & ~n501;
  assign n6687 = ~n1027 & ~n1145;
  assign n6688 = n6686 & n6687;
  assign n6689 = n6685 & n6688;
  assign n6690 = ~n2335 & ~n2664;
  assign n6691 = n4798 & n6690;
  assign n6692 = n4790 & n6691;
  assign n6693 = n6689 & n6692;
  assign n6694 = n6683 & n6693;
  assign n6695 = ~n1172 & n6694;
  assign n6696 = ~n1054 & n6695;
  assign n6697 = ~n996 & n6696;
  assign n6698 = ~n2306 & ~n2362;
  assign n6699 = n6697 & n6698;
  assign n6700 = n6677 & n6699;
  assign n6701 = ~n4549 & ~n4647;
  assign n6702 = ~n5497 & ~n5555;
  assign n6703 = n6701 & n6702;
  assign n6704 = ~n2691 & ~n3552;
  assign n6705 = ~n3254 & ~n4766;
  assign n6706 = n6704 & n6705;
  assign n6707 = n6703 & n6706;
  assign n6708 = n6700 & n6707;
  assign n6709 = ~n2049 & ~n2080;
  assign n6710 = n3808 & n6709;
  assign n6711 = n3823 & n6710;
  assign n6712 = n6708 & n6711;
  assign n6713 = n6676 & n6712;
  assign n6714 = n6284 & n6713;
  assign n6715 = ~n6195 & ~n6714;
  assign n6716 = ~n6120 & n6715;
  assign po007 = n6115 | ~n6716;
  assign n6718 = n5886 & ~n5943;
  assign n6719 = n5859 & ~n6001;
  assign n6720 = ~n5827 & n5885;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n6718 & n6721;
  assign n6723 = ~n1115 & ~n1144;
  assign n6724 = n1056 & n6723;
  assign n6725 = ~n1208 & n6724;
  assign n6726 = n4920 & n6725;
  assign n6727 = n5873 & n6726;
  assign n6728 = n4932 & n6727;
  assign n6729 = ~n5865 & n6728;
  assign n6730 = ~n1372 & n6729;
  assign n6731 = ~n2243 & n6730;
  assign n6732 = ~n3104 & n6731;
  assign n6733 = ~n3971 & n6732;
  assign n6734 = ~n4003 & n6733;
  assign n6735 = ~n4872 & n6734;
  assign n6736 = ~n5801 & n6735;
  assign n6737 = ~n5864 & n6736;
  assign n6738 = n5891 & n6737;
  assign n6739 = n5863 & n6738;
  assign n6740 = ~n5528 & ~n6144;
  assign n6741 = n5757 & n6740;
  assign n6742 = n5759 & n6741;
  assign n6743 = n5756 & n6742;
  assign n6744 = n5753 & n6743;
  assign n6745 = ~n1172 & n6744;
  assign n6746 = ~n996 & n6745;
  assign n6747 = ~n2306 & n6746;
  assign n6748 = n3819 & n6747;
  assign n6749 = n3821 & n6748;
  assign n6750 = n6183 & n6749;
  assign n6751 = n5741 & n6750;
  assign n6752 = ~n6137 & n6751;
  assign n6753 = n6193 & n6752;
  assign n6754 = n6134 & n6753;
  assign n6755 = n1357 & ~n6754;
  assign n6756 = n5888 & ~n6027;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = ~n6739 & n6757;
  assign n6759 = n5889 & ~n6056;
  assign n6760 = n5860 & ~n5967;
  assign n6761 = n5864 & ~n5917;
  assign n6762 = ~n2694 & ~n3227;
  assign n6763 = n6678 & n6762;
  assign n6764 = ~n3256 & ~n3525;
  assign n6765 = n3941 & n6764;
  assign n6766 = n6763 & n6765;
  assign n6767 = n5758 & n6766;
  assign n6768 = ~n1027 & ~n2021;
  assign n6769 = n3858 & n6768;
  assign n6770 = n2246 & n5713;
  assign n6771 = n6769 & n6770;
  assign n6772 = n3859 & n6690;
  assign n6773 = n5718 & n6772;
  assign n6774 = n6771 & n6773;
  assign n6775 = n6767 & n6774;
  assign n6776 = ~n1172 & n6775;
  assign n6777 = ~n1054 & n6776;
  assign n6778 = ~n996 & n6777;
  assign n6779 = n6698 & n6778;
  assign n6780 = n6677 & n6779;
  assign n6781 = n6707 & n6780;
  assign n6782 = n6711 & n6781;
  assign n6783 = n6676 & n6782;
  assign n6784 = n6284 & n6783;
  assign n6785 = n1055 & ~n6784;
  assign n6786 = ~n1026 & n5867;
  assign n6787 = ~n1086 & ~n1299;
  assign n6788 = n6786 & n6787;
  assign n6789 = n1239 & n6788;
  assign n6790 = ~n1270 & n6789;
  assign n6791 = n844 & n6790;
  assign n6792 = ~n1372 & n6791;
  assign n6793 = ~n2243 & n6792;
  assign n6794 = ~n6785 & n6793;
  assign n6795 = ~n3104 & n6794;
  assign n6796 = ~n3971 & n6795;
  assign n6797 = ~n4003 & n6796;
  assign n6798 = ~n4872 & n6797;
  assign n6799 = ~n5801 & n6798;
  assign n6800 = ~n6761 & n6799;
  assign n6801 = ~n6760 & n6800;
  assign n6802 = ~n6759 & n6801;
  assign n6803 = n5865 & ~n6114;
  assign n6804 = ~n1804 & n3082;
  assign n6805 = ~n1649 & ~n2050;
  assign n6806 = n3085 & n6805;
  assign n6807 = n3089 & n6806;
  assign n6808 = n4954 & n4955;
  assign n6809 = n6807 & n6808;
  assign n6810 = n6804 & n6809;
  assign n6811 = ~n5834 & n6810;
  assign n6812 = ~n2242 & n6811;
  assign n6813 = ~n3095 & n6812;
  assign n6814 = ~n3997 & n6813;
  assign n6815 = ~n4003 & n6814;
  assign n6816 = ~n4837 & n6815;
  assign n6817 = ~n5822 & n6816;
  assign n6818 = ~n5833 & n6817;
  assign n6819 = n5856 & n6818;
  assign n6820 = n5832 & n6819;
  assign n6821 = n5861 & ~n6820;
  assign n6822 = ~n6803 & ~n6821;
  assign n6823 = n6802 & n6822;
  assign n6824 = n6758 & n6823;
  assign n6825 = n6722 & n6824;
  assign n6826 = n5830 & ~n6739;
  assign n6827 = ~n5827 & n5850;
  assign n6828 = n5828 & ~n6001;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = ~n6826 & n6829;
  assign n6831 = n5853 & ~n6027;
  assign n6832 = n5829 & ~n5967;
  assign n6833 = n1927 & ~n6754;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = ~n6831 & n6834;
  assign n6836 = n5851 & ~n5943;
  assign n6837 = n5833 & ~n5917;
  assign n6838 = n2050 & ~n6784;
  assign n6839 = n3889 & n5835;
  assign n6840 = ~n1649 & ~n2020;
  assign n6841 = n2207 & n6840;
  assign n6842 = n4955 & n6841;
  assign n6843 = n4954 & n6842;
  assign n6844 = n6839 & n6843;
  assign n6845 = ~n6838 & n6844;
  assign n6846 = ~n2242 & n6845;
  assign n6847 = ~n3095 & n6846;
  assign n6848 = ~n3997 & n6847;
  assign n6849 = ~n4003 & n6848;
  assign n6850 = ~n4837 & n6849;
  assign n6851 = ~n5822 & n6850;
  assign n6852 = ~n6837 & n6851;
  assign n6853 = ~n6820 & n6852;
  assign n6854 = ~n6836 & n6853;
  assign n6855 = n5854 & ~n6056;
  assign n6856 = n5834 & ~n6114;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = n6854 & n6857;
  assign n6859 = n6835 & n6858;
  assign n6860 = n6830 & n6859;
  assign n6861 = ~n6825 & ~n6860;
  assign n6862 = n5748 & ~n5943;
  assign n6863 = n5786 & ~n6001;
  assign n6864 = n5823 & ~n6820;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = ~n6862 & n6865;
  assign n6867 = n5746 & ~n6027;
  assign n6868 = n5747 & ~n5967;
  assign n6869 = n2965 & ~n6754;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = ~n6867 & n6870;
  assign n6872 = n5809 & ~n6056;
  assign n6873 = n5751 & ~n5917;
  assign n6874 = n2363 & ~n6784;
  assign n6875 = ~n2934 & n3054;
  assign n6876 = n2573 & n5002;
  assign n6877 = n5897 & n6876;
  assign n6878 = n6875 & n6877;
  assign n6879 = ~n6874 & n6878;
  assign n6880 = ~n3066 & n6879;
  assign n6881 = ~n3983 & n6880;
  assign n6882 = ~n4003 & n6881;
  assign n6883 = ~n4024 & n6882;
  assign n6884 = ~n4999 & n6883;
  assign n6885 = ~n6873 & n6884;
  assign n6886 = ~n5827 & n6885;
  assign n6887 = ~n6872 & n6886;
  assign n6888 = n5770 & ~n6114;
  assign n6889 = n5802 & ~n6739;
  assign n6890 = ~n6888 & ~n6889;
  assign n6891 = n6887 & n6890;
  assign n6892 = n6871 & n6891;
  assign n6893 = n6866 & n6892;
  assign n6894 = ~n6861 & ~n6893;
  assign n6895 = pi005 & ~n2543;
  assign n6896 = n5772 & n6895;
  assign n6897 = n5776 & n6896;
  assign n6898 = n6875 & n6897;
  assign n6899 = ~n6874 & n6898;
  assign n6900 = ~n3066 & n6899;
  assign n6901 = ~n3983 & n6900;
  assign n6902 = ~n4003 & n6901;
  assign n6903 = ~n4024 & n6902;
  assign n6904 = ~n4999 & n6903;
  assign n6905 = ~n6873 & n6904;
  assign n6906 = ~n5827 & n6905;
  assign n6907 = ~n6872 & n6906;
  assign n6908 = n6890 & n6907;
  assign n6909 = n6871 & n6908;
  assign n6910 = n6866 & n6909;
  assign n6911 = n5914 & ~n6820;
  assign n6912 = n5912 & ~n5917;
  assign n6913 = ~n6911 & n6912;
  assign n6914 = ~n5827 & n5909;
  assign n6915 = n5915 & ~n6739;
  assign n6916 = ~n6914 & ~n6915;
  assign n6917 = n6913 & n6916;
  assign n6918 = ~n6910 & ~n6917;
  assign n6919 = ~n6894 & n6918;
  assign n6920 = ~n5827 & n5938;
  assign n6921 = n5920 & ~n6820;
  assign n6922 = n5918 & ~n6739;
  assign n6923 = ~n6921 & ~n6922;
  assign n6924 = ~n6920 & n6923;
  assign n6925 = n5935 & ~n5967;
  assign n6926 = n5936 & ~n6027;
  assign n6927 = n3493 & ~n6754;
  assign n6928 = ~n6926 & ~n6927;
  assign n6929 = ~n6925 & n6928;
  assign n6930 = n5919 & ~n6001;
  assign n6931 = ~n5917 & n5923;
  assign n6932 = n3553 & ~n6784;
  assign n6933 = ~n3136 & ~n3464;
  assign n6934 = ~n3165 & n6933;
  assign n6935 = ~n3524 & ~n3710;
  assign n6936 = n5062 & n6935;
  assign n6937 = n5948 & n6936;
  assign n6938 = n6934 & n6937;
  assign n6939 = ~n6932 & n6938;
  assign n6940 = ~n3940 & n6939;
  assign n6941 = ~n4001 & n6940;
  assign n6942 = ~n5043 & n6941;
  assign n6943 = ~n6931 & n6942;
  assign n6944 = ~n5943 & n6943;
  assign n6945 = ~n6930 & n6944;
  assign n6946 = n5939 & ~n6056;
  assign n6947 = n5924 & ~n6114;
  assign n6948 = ~n6946 & ~n6947;
  assign n6949 = n6945 & n6948;
  assign n6950 = n6929 & n6949;
  assign n6951 = n6924 & n6950;
  assign n6952 = n5047 & ~n5911;
  assign n6953 = ~n5917 & n6952;
  assign n6954 = ~n6911 & n6953;
  assign n6955 = n6916 & n6954;
  assign n6956 = ~n6951 & ~n6955;
  assign n6957 = ~n6919 & n6956;
  assign n6958 = ~n5943 & n5963;
  assign n6959 = n5958 & ~n5967;
  assign n6960 = ~n6931 & n6959;
  assign n6961 = ~n6958 & n6960;
  assign n6962 = ~n5827 & n5964;
  assign n6963 = n5960 & ~n6820;
  assign n6964 = n5961 & ~n6739;
  assign n6965 = ~n6963 & ~n6964;
  assign n6966 = ~n6962 & n6965;
  assign n6967 = n6961 & n6966;
  assign n6968 = n3800 & n4094;
  assign n6969 = n5927 & n6968;
  assign n6970 = n6934 & n6969;
  assign n6971 = ~n6932 & n6970;
  assign n6972 = ~n3940 & n6971;
  assign n6973 = ~n4001 & n6972;
  assign n6974 = ~n5043 & n6973;
  assign n6975 = ~n6931 & n6974;
  assign n6976 = ~n5943 & n6975;
  assign n6977 = ~n6930 & n6976;
  assign n6978 = n6948 & n6977;
  assign n6979 = n6929 & n6978;
  assign n6980 = n6924 & n6979;
  assign n6981 = ~n6967 & ~n6980;
  assign n6982 = ~n6957 & n6981;
  assign n6983 = ~n5967 & n5977;
  assign n6984 = ~n6931 & n6983;
  assign n6985 = ~n6958 & n6984;
  assign n6986 = n6966 & n6985;
  assign n6987 = ~n5943 & n5997;
  assign n6988 = n5985 & ~n6114;
  assign n6989 = n5996 & ~n6056;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = ~n6987 & n6990;
  assign n6992 = n5981 & ~n6027;
  assign n6993 = n4222 & ~n6754;
  assign n6994 = ~n6959 & ~n6993;
  assign n6995 = ~n6992 & n6994;
  assign n6996 = n5982 & ~n6820;
  assign n6997 = n4550 & ~n6784;
  assign n6998 = ~n4192 & n4892;
  assign n6999 = ~n4608 & n5090;
  assign n7000 = n5095 & n6999;
  assign n7001 = n5987 & n7000;
  assign n7002 = n6998 & n7001;
  assign n7003 = ~n6997 & n7002;
  assign n7004 = ~n4817 & n7003;
  assign n7005 = ~n4902 & n7004;
  assign n7006 = ~n6931 & n7005;
  assign n7007 = ~n6001 & n7006;
  assign n7008 = ~n6996 & n7007;
  assign n7009 = n5980 & ~n6739;
  assign n7010 = ~n5827 & n5994;
  assign n7011 = ~n7009 & ~n7010;
  assign n7012 = n7008 & n7011;
  assign n7013 = n6995 & n7012;
  assign n7014 = n6991 & n7013;
  assign n7015 = ~n6986 & ~n7014;
  assign n7016 = ~n6982 & n7015;
  assign n7017 = ~n6001 & n6016;
  assign n7018 = n6019 & ~n6820;
  assign n7019 = ~n5943 & n6018;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = ~n7017 & n7020;
  assign n7022 = n6022 & ~n6027;
  assign n7023 = ~n6931 & n7022;
  assign n7024 = ~n6959 & n7023;
  assign n7025 = ~n5827 & n6024;
  assign n7026 = n6015 & ~n6739;
  assign n7027 = ~n7025 & ~n7026;
  assign n7028 = n7024 & n7027;
  assign n7029 = n7021 & n7028;
  assign n7030 = n4431 & n4737;
  assign n7031 = n6004 & n7030;
  assign n7032 = n4371 & n4609;
  assign n7033 = n4312 & n4490;
  assign n7034 = n7032 & n7033;
  assign n7035 = n7031 & n7034;
  assign n7036 = n6998 & n7035;
  assign n7037 = ~n6997 & n7036;
  assign n7038 = ~n4817 & n7037;
  assign n7039 = ~n4902 & n7038;
  assign n7040 = ~n6931 & n7039;
  assign n7041 = ~n6001 & n7040;
  assign n7042 = ~n6996 & n7041;
  assign n7043 = n7011 & n7042;
  assign n7044 = n6995 & n7043;
  assign n7045 = n6991 & n7044;
  assign n7046 = ~n7029 & ~n7045;
  assign n7047 = ~n7016 & n7046;
  assign n7048 = ~n5943 & n6051;
  assign n7049 = n6035 & ~n6114;
  assign n7050 = n6032 & ~n6820;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = ~n7048 & n7051;
  assign n7053 = n5141 & ~n6754;
  assign n7054 = ~n6959 & ~n7022;
  assign n7055 = ~n7053 & n7054;
  assign n7056 = ~n5827 & n6031;
  assign n7057 = n5498 & ~n6784;
  assign n7058 = ~n5199 & n6036;
  assign n7059 = n5319 & ~n5527;
  assign n7060 = n6043 & n7059;
  assign n7061 = n6040 & n7060;
  assign n7062 = n7058 & n7061;
  assign n7063 = ~n7057 & n7062;
  assign n7064 = ~n5808 & n7063;
  assign n7065 = ~n6931 & n7064;
  assign n7066 = ~n6056 & n7065;
  assign n7067 = ~n7056 & n7066;
  assign n7068 = ~n6001 & n6052;
  assign n7069 = n6030 & ~n6739;
  assign n7070 = ~n7068 & ~n7069;
  assign n7071 = n7067 & n7070;
  assign n7072 = n7055 & n7071;
  assign n7073 = n7052 & n7072;
  assign n7074 = ~n6027 & n6058;
  assign n7075 = ~n6931 & n7074;
  assign n7076 = ~n6959 & n7075;
  assign n7077 = n7027 & n7076;
  assign n7078 = n7021 & n7077;
  assign n7079 = ~n7073 & ~n7078;
  assign n7080 = ~n7047 & n7079;
  assign n7081 = ~n6056 & n6093;
  assign n7082 = ~n5943 & n6110;
  assign n7083 = ~n7081 & ~n7082;
  assign n7084 = ~n6001 & n6092;
  assign n7085 = ~n5827 & n6101;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = n7083 & n7086;
  assign n7088 = ~n5769 & ~n6931;
  assign n7089 = ~n6114 & n7088;
  assign n7090 = n7054 & n7089;
  assign n7091 = n6107 & ~n6820;
  assign n7092 = n6090 & ~n6739;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = n7090 & n7093;
  assign n7095 = n7087 & n7094;
  assign n7096 = n6064 & n6068;
  assign n7097 = n6067 & n7096;
  assign n7098 = n6071 & n6074;
  assign n7099 = n6065 & n6073;
  assign n7100 = n7098 & n7099;
  assign n7101 = n7097 & n7100;
  assign n7102 = n7058 & n7101;
  assign n7103 = ~n7057 & n7102;
  assign n7104 = ~n5808 & n7103;
  assign n7105 = ~n6931 & n7104;
  assign n7106 = ~n6056 & n7105;
  assign n7107 = ~n7056 & n7106;
  assign n7108 = n7070 & n7107;
  assign n7109 = n7055 & n7108;
  assign n7110 = n7052 & n7109;
  assign n7111 = ~n7095 & ~n7110;
  assign n7112 = ~n7080 & n7111;
  assign n7113 = ~n2050 & ~n2242;
  assign n7114 = ~n3095 & n7113;
  assign n7115 = ~n3997 & n7114;
  assign n7116 = ~n4837 & n7115;
  assign n7117 = ~n5822 & n7116;
  assign n7118 = ~n6820 & n7117;
  assign n7119 = ~n1055 & ~n1372;
  assign n7120 = ~n2243 & n7119;
  assign n7121 = ~n3104 & n7120;
  assign n7122 = ~n3971 & n7121;
  assign n7123 = ~n4872 & n7122;
  assign n7124 = ~n5801 & n7123;
  assign n7125 = ~n6739 & n7124;
  assign n7126 = ~n2363 & ~n3066;
  assign n7127 = ~n3983 & n7126;
  assign n7128 = ~n4024 & n7127;
  assign n7129 = ~n4999 & n7128;
  assign n7130 = ~n5827 & n7129;
  assign n7131 = ~n7125 & ~n7130;
  assign n7132 = ~n7118 & n7131;
  assign n7133 = n6403 & n6462;
  assign n7134 = n6523 & ~n6552;
  assign n7135 = n6674 & n7134;
  assign n7136 = n7133 & n7135;
  assign n7137 = n6284 & n7136;
  assign n7138 = ~n6784 & n7137;
  assign n7139 = ~n6931 & n7138;
  assign n7140 = ~n6959 & n7139;
  assign n7141 = n6553 & ~n6754;
  assign n7142 = ~n7022 & ~n7141;
  assign n7143 = n7140 & n7142;
  assign n7144 = ~n4550 & ~n4817;
  assign n7145 = ~n4902 & n7144;
  assign n7146 = ~n6001 & n7145;
  assign n7147 = ~n3553 & ~n3940;
  assign n7148 = ~n4001 & n7147;
  assign n7149 = ~n5043 & n7148;
  assign n7150 = ~n5943 & n7149;
  assign n7151 = ~n7146 & ~n7150;
  assign n7152 = ~n5769 & ~n6114;
  assign n7153 = ~n5498 & ~n5808;
  assign n7154 = ~n6056 & n7153;
  assign n7155 = ~n7152 & ~n7154;
  assign n7156 = n7151 & n7155;
  assign n7157 = n7143 & n7156;
  assign n7158 = n7132 & n7157;
  assign n7159 = ~pi012 & ~n5769;
  assign n7160 = ~n6931 & n7159;
  assign n7161 = ~n6114 & n7160;
  assign n7162 = n7054 & n7161;
  assign n7163 = n7093 & n7162;
  assign n7164 = n7087 & n7163;
  assign n7165 = ~n7158 & ~n7164;
  assign n7166 = ~n7112 & n7165;
  assign n7167 = pi013 & ~n6432;
  assign n7168 = ~n6313 & ~n6461;
  assign n7169 = ~n6342 & ~n6372;
  assign n7170 = n7168 & n7169;
  assign n7171 = n7167 & n7170;
  assign n7172 = ~n6493 & ~n6672;
  assign n7173 = ~n6522 & ~n6552;
  assign n7174 = n7172 & n7173;
  assign n7175 = ~n6401 & ~n6584;
  assign n7176 = ~n6613 & ~n6643;
  assign n7177 = n7175 & n7176;
  assign n7178 = n7174 & n7177;
  assign n7179 = n7171 & n7178;
  assign n7180 = n6284 & n7179;
  assign n7181 = ~n6784 & n7180;
  assign n7182 = ~n6931 & n7181;
  assign n7183 = ~n6959 & n7182;
  assign n7184 = n7142 & n7183;
  assign n7185 = n7156 & n7184;
  assign n7186 = n7132 & n7185;
  assign n7187 = ~n7166 & ~n7186;
  assign n7188 = ~n5943 & n6137;
  assign n7189 = n6125 & ~n6820;
  assign n7190 = ~n6056 & n6132;
  assign n7191 = ~n7189 & ~n7190;
  assign n7192 = ~n7188 & n7191;
  assign n7193 = ~n6553 & ~n6784;
  assign n7194 = ~n6754 & ~n7193;
  assign n7195 = ~n6931 & n7194;
  assign n7196 = n7054 & n7195;
  assign n7197 = ~n5827 & n6192;
  assign n7198 = ~n7152 & ~n7197;
  assign n7199 = ~n6001 & n6188;
  assign n7200 = n6131 & ~n6739;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = n7198 & n7201;
  assign n7203 = n7196 & n7202;
  assign n7204 = n7192 & n7203;
  assign n7205 = ~n7187 & ~n7204;
  assign n7206 = pi014 & ~n7193;
  assign n7207 = ~n6754 & n7206;
  assign n7208 = ~n6931 & n7207;
  assign n7209 = n7054 & n7208;
  assign n7210 = n7202 & n7209;
  assign n7211 = n7192 & n7210;
  assign n7212 = ~n1299 & ~n1372;
  assign n7213 = ~n2243 & n7212;
  assign n7214 = ~n3104 & n7213;
  assign n7215 = ~n3971 & n7214;
  assign n7216 = ~n4872 & n7215;
  assign n7217 = ~n5801 & n7216;
  assign n7218 = ~n6739 & n7217;
  assign n7219 = ~n3053 & ~n3066;
  assign n7220 = ~n3983 & n7219;
  assign n7221 = ~n4024 & n7220;
  assign n7222 = ~n4999 & n7221;
  assign n7223 = ~n5827 & n7222;
  assign n7224 = ~n1804 & ~n2242;
  assign n7225 = ~n3095 & n7224;
  assign n7226 = ~n3997 & n7225;
  assign n7227 = ~n4837 & n7226;
  assign n7228 = ~n5822 & n7227;
  assign n7229 = ~n6820 & n7228;
  assign n7230 = ~n7223 & ~n7229;
  assign n7231 = ~n7218 & n7230;
  assign n7232 = ~n3136 & ~n3940;
  assign n7233 = ~n4001 & n7232;
  assign n7234 = ~n5043 & n7233;
  assign n7235 = ~n5943 & n7234;
  assign n7236 = ~n6253 & ~n6784;
  assign n7237 = pi016 & ~n501;
  assign n7238 = n5713 & n7237;
  assign n7239 = n6138 & n7238;
  assign n7240 = ~pi151 & pi159;
  assign n7241 = ~n6144 & ~n7240;
  assign n7242 = n5720 & n7241;
  assign n7243 = n4797 & n7242;
  assign n7244 = n6143 & n7243;
  assign n7245 = n7239 & n7244;
  assign n7246 = ~n1172 & n7245;
  assign n7247 = ~n996 & n7246;
  assign n7248 = ~n2306 & n7247;
  assign n7249 = ~n500 & n7248;
  assign n7250 = n6677 & n7249;
  assign n7251 = pi153 & ~pi161;
  assign n7252 = ~pi154 & pi162;
  assign n7253 = pi154 & ~pi162;
  assign n7254 = ~pi155 & pi163;
  assign n7255 = pi155 & ~pi163;
  assign n7256 = ~pi156 & pi164;
  assign n7257 = pi156 & ~pi164;
  assign n7258 = pi158 & ~pi166;
  assign n7259 = pi157 & ~pi165;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = ~pi157 & pi165;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7257 & ~n7262;
  assign n7264 = ~n7256 & ~n7263;
  assign n7265 = ~n7255 & ~n7264;
  assign n7266 = ~n7254 & ~n7265;
  assign n7267 = ~n7253 & ~n7266;
  assign n7268 = ~n7252 & ~n7267;
  assign n7269 = ~n7251 & ~n7268;
  assign n7270 = ~pi153 & pi161;
  assign n7271 = ~pi152 & pi160;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = ~n7269 & n7272;
  assign n7274 = pi151 & ~pi159;
  assign n7275 = pi152 & ~pi160;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = ~n7273 & n7276;
  assign n7278 = n6181 & ~n7277;
  assign n7279 = n4788 & n5732;
  assign n7280 = n7278 & n7279;
  assign n7281 = n7250 & n7280;
  assign n7282 = ~n562 & ~n2080;
  assign n7283 = n2316 & n7282;
  assign n7284 = n4787 & n7283;
  assign n7285 = n7281 & n7284;
  assign n7286 = ~n7236 & n7285;
  assign n7287 = ~n6137 & n7286;
  assign n7288 = n6193 & n7287;
  assign n7289 = n6134 & n7288;
  assign n7290 = ~n7235 & n7289;
  assign n7291 = ~n4521 & ~n4817;
  assign n7292 = ~n4902 & n7291;
  assign n7293 = ~n6001 & n7292;
  assign n7294 = ~n5199 & ~n5808;
  assign n7295 = ~n6056 & n7294;
  assign n7296 = ~n7293 & ~n7295;
  assign n7297 = n7290 & n7296;
  assign n7298 = n7231 & n7297;
  assign n7299 = ~pi151 & pi183;
  assign n7300 = pi153 & ~pi185;
  assign n7301 = ~pi154 & pi186;
  assign n7302 = pi154 & ~pi186;
  assign n7303 = ~pi155 & pi187;
  assign n7304 = pi155 & ~pi187;
  assign n7305 = ~pi156 & pi188;
  assign n7306 = pi156 & ~pi188;
  assign n7307 = pi158 & ~pi190;
  assign n7308 = pi157 & ~pi189;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~pi157 & pi189;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~n7306 & ~n7311;
  assign n7313 = ~n7305 & ~n7312;
  assign n7314 = ~n7304 & ~n7313;
  assign n7315 = ~n7303 & ~n7314;
  assign n7316 = ~n7302 & ~n7315;
  assign n7317 = ~n7301 & ~n7316;
  assign n7318 = ~n7300 & ~n7317;
  assign n7319 = ~pi153 & pi185;
  assign n7320 = ~pi152 & pi184;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = ~n7318 & n7321;
  assign n7323 = pi151 & ~pi183;
  assign n7324 = pi152 & ~pi184;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~n7322 & n7325;
  assign n7327 = ~n7299 & ~n7326;
  assign n7328 = ~pi151 & pi223;
  assign n7329 = pi153 & ~pi225;
  assign n7330 = ~pi154 & pi226;
  assign n7331 = pi154 & ~pi226;
  assign n7332 = ~pi155 & pi227;
  assign n7333 = pi155 & ~pi227;
  assign n7334 = ~pi156 & pi228;
  assign n7335 = pi156 & ~pi228;
  assign n7336 = pi158 & ~pi230;
  assign n7337 = pi157 & ~pi229;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~pi157 & pi229;
  assign n7340 = ~n7338 & ~n7339;
  assign n7341 = ~n7335 & ~n7340;
  assign n7342 = ~n7334 & ~n7341;
  assign n7343 = ~n7333 & ~n7342;
  assign n7344 = ~n7332 & ~n7343;
  assign n7345 = ~n7331 & ~n7344;
  assign n7346 = ~n7330 & ~n7345;
  assign n7347 = ~n7329 & ~n7346;
  assign n7348 = ~pi153 & pi225;
  assign n7349 = ~pi152 & pi224;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = ~n7347 & n7350;
  assign n7352 = pi151 & ~pi223;
  assign n7353 = pi152 & ~pi224;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n7351 & n7354;
  assign n7356 = ~n7328 & ~n7355;
  assign n7357 = ~n7327 & ~n7356;
  assign n7358 = ~pi151 & pi199;
  assign n7359 = pi153 & ~pi201;
  assign n7360 = ~pi154 & pi202;
  assign n7361 = pi154 & ~pi202;
  assign n7362 = ~pi155 & pi203;
  assign n7363 = pi155 & ~pi203;
  assign n7364 = ~pi156 & pi204;
  assign n7365 = pi156 & ~pi204;
  assign n7366 = pi158 & ~pi206;
  assign n7367 = pi157 & ~pi205;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~pi157 & pi205;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n7365 & ~n7370;
  assign n7372 = ~n7364 & ~n7371;
  assign n7373 = ~n7363 & ~n7372;
  assign n7374 = ~n7362 & ~n7373;
  assign n7375 = ~n7361 & ~n7374;
  assign n7376 = ~n7360 & ~n7375;
  assign n7377 = ~n7359 & ~n7376;
  assign n7378 = ~pi153 & pi201;
  assign n7379 = ~pi152 & pi200;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = ~n7377 & n7380;
  assign n7382 = pi151 & ~pi199;
  assign n7383 = pi152 & ~pi200;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = ~n7381 & n7384;
  assign n7386 = ~n7358 & ~n7385;
  assign n7387 = ~pi151 & pi207;
  assign n7388 = pi153 & ~pi209;
  assign n7389 = ~pi154 & pi210;
  assign n7390 = pi154 & ~pi210;
  assign n7391 = ~pi155 & pi211;
  assign n7392 = pi155 & ~pi211;
  assign n7393 = ~pi156 & pi212;
  assign n7394 = pi156 & ~pi212;
  assign n7395 = pi158 & ~pi214;
  assign n7396 = pi157 & ~pi213;
  assign n7397 = ~n7395 & ~n7396;
  assign n7398 = ~pi157 & pi213;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = ~n7394 & ~n7399;
  assign n7401 = ~n7393 & ~n7400;
  assign n7402 = ~n7392 & ~n7401;
  assign n7403 = ~n7391 & ~n7402;
  assign n7404 = ~n7390 & ~n7403;
  assign n7405 = ~n7389 & ~n7404;
  assign n7406 = ~n7388 & ~n7405;
  assign n7407 = ~pi153 & pi209;
  assign n7408 = ~pi152 & pi208;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = ~n7406 & n7409;
  assign n7411 = pi151 & ~pi207;
  assign n7412 = pi152 & ~pi208;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = ~n7410 & n7413;
  assign n7415 = ~n7387 & ~n7414;
  assign n7416 = ~n7386 & ~n7415;
  assign n7417 = n7357 & n7416;
  assign n7418 = ~pi151 & pi215;
  assign n7419 = pi153 & ~pi217;
  assign n7420 = ~pi154 & pi218;
  assign n7421 = pi154 & ~pi218;
  assign n7422 = ~pi155 & pi219;
  assign n7423 = pi155 & ~pi219;
  assign n7424 = ~pi156 & pi220;
  assign n7425 = pi156 & ~pi220;
  assign n7426 = pi158 & ~pi222;
  assign n7427 = pi157 & ~pi221;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = ~pi157 & pi221;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~n7425 & ~n7430;
  assign n7432 = ~n7424 & ~n7431;
  assign n7433 = ~n7423 & ~n7432;
  assign n7434 = ~n7422 & ~n7433;
  assign n7435 = ~n7421 & ~n7434;
  assign n7436 = ~n7420 & ~n7435;
  assign n7437 = ~n7419 & ~n7436;
  assign n7438 = ~pi153 & pi217;
  assign n7439 = ~pi152 & pi216;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = ~n7437 & n7440;
  assign n7442 = pi151 & ~pi215;
  assign n7443 = pi152 & ~pi216;
  assign n7444 = ~n7442 & ~n7443;
  assign n7445 = ~n7441 & n7444;
  assign n7446 = ~n7418 & ~n7445;
  assign n7447 = ~pi151 & pi247;
  assign n7448 = pi153 & ~pi249;
  assign n7449 = ~pi154 & pi250;
  assign n7450 = pi154 & ~pi250;
  assign n7451 = ~pi155 & pi251;
  assign n7452 = pi155 & ~pi251;
  assign n7453 = ~pi156 & pi252;
  assign n7454 = pi156 & ~pi252;
  assign n7455 = pi158 & ~pi254;
  assign n7456 = pi157 & ~pi253;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~pi157 & pi253;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = ~n7454 & ~n7459;
  assign n7461 = ~n7453 & ~n7460;
  assign n7462 = ~n7452 & ~n7461;
  assign n7463 = ~n7451 & ~n7462;
  assign n7464 = ~n7450 & ~n7463;
  assign n7465 = ~n7449 & ~n7464;
  assign n7466 = ~n7448 & ~n7465;
  assign n7467 = ~pi153 & pi249;
  assign n7468 = ~pi152 & pi248;
  assign n7469 = ~n7467 & ~n7468;
  assign n7470 = ~n7466 & n7469;
  assign n7471 = pi151 & ~pi247;
  assign n7472 = pi152 & ~pi248;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = ~n7470 & n7473;
  assign n7475 = ~n7447 & ~n7474;
  assign n7476 = ~n7446 & ~n7475;
  assign n7477 = ~pi151 & pi263;
  assign n7478 = pi153 & ~pi265;
  assign n7479 = ~pi154 & pi266;
  assign n7480 = pi154 & ~pi266;
  assign n7481 = ~pi155 & pi267;
  assign n7482 = pi155 & ~pi267;
  assign n7483 = ~pi156 & pi268;
  assign n7484 = pi156 & ~pi268;
  assign n7485 = pi158 & ~pi270;
  assign n7486 = pi157 & ~pi269;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = ~pi157 & pi269;
  assign n7489 = ~n7487 & ~n7488;
  assign n7490 = ~n7484 & ~n7489;
  assign n7491 = ~n7483 & ~n7490;
  assign n7492 = ~n7482 & ~n7491;
  assign n7493 = ~n7481 & ~n7492;
  assign n7494 = ~n7480 & ~n7493;
  assign n7495 = ~n7479 & ~n7494;
  assign n7496 = ~n7478 & ~n7495;
  assign n7497 = ~pi153 & pi265;
  assign n7498 = ~pi152 & pi264;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = ~n7496 & n7499;
  assign n7501 = pi151 & ~pi263;
  assign n7502 = pi152 & ~pi264;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = ~n7500 & n7503;
  assign n7505 = ~n7477 & ~n7504;
  assign n7506 = ~pi151 & pi167;
  assign n7507 = pi153 & ~pi169;
  assign n7508 = ~pi154 & pi170;
  assign n7509 = pi154 & ~pi170;
  assign n7510 = ~pi155 & pi171;
  assign n7511 = pi155 & ~pi171;
  assign n7512 = ~pi156 & pi172;
  assign n7513 = pi156 & ~pi172;
  assign n7514 = pi158 & ~pi174;
  assign n7515 = pi157 & ~pi173;
  assign n7516 = ~n7514 & ~n7515;
  assign n7517 = ~pi157 & pi173;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~n7513 & ~n7518;
  assign n7520 = ~n7512 & ~n7519;
  assign n7521 = ~n7511 & ~n7520;
  assign n7522 = ~n7510 & ~n7521;
  assign n7523 = ~n7509 & ~n7522;
  assign n7524 = ~n7508 & ~n7523;
  assign n7525 = ~n7507 & ~n7524;
  assign n7526 = ~pi153 & pi169;
  assign n7527 = ~pi152 & pi168;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = ~n7525 & n7528;
  assign n7530 = pi151 & ~pi167;
  assign n7531 = pi152 & ~pi168;
  assign n7532 = ~n7530 & ~n7531;
  assign n7533 = ~n7529 & n7532;
  assign n7534 = ~n7506 & ~n7533;
  assign n7535 = ~n7505 & ~n7534;
  assign n7536 = n7476 & n7535;
  assign n7537 = n7417 & n7536;
  assign n7538 = ~pi151 & pi175;
  assign n7539 = pi151 & ~pi175;
  assign n7540 = ~pi152 & pi176;
  assign n7541 = pi152 & ~pi176;
  assign n7542 = ~pi153 & pi177;
  assign n7543 = pi153 & ~pi177;
  assign n7544 = ~pi154 & pi178;
  assign n7545 = pi154 & ~pi178;
  assign n7546 = ~pi155 & pi179;
  assign n7547 = pi155 & ~pi179;
  assign n7548 = ~pi156 & pi180;
  assign n7549 = pi156 & ~pi180;
  assign n7550 = pi158 & ~pi182;
  assign n7551 = pi157 & ~pi181;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = ~pi157 & pi181;
  assign n7554 = ~n7552 & ~n7553;
  assign n7555 = ~n7549 & ~n7554;
  assign n7556 = ~n7548 & ~n7555;
  assign n7557 = ~n7547 & ~n7556;
  assign n7558 = ~n7546 & ~n7557;
  assign n7559 = ~n7545 & ~n7558;
  assign n7560 = ~n7544 & ~n7559;
  assign n7561 = ~n7543 & ~n7560;
  assign n7562 = ~n7542 & ~n7561;
  assign n7563 = ~n7541 & ~n7562;
  assign n7564 = ~n7540 & ~n7563;
  assign n7565 = ~n7539 & ~n7564;
  assign n7566 = ~n7538 & ~n7565;
  assign n7567 = ~pi151 & pi191;
  assign n7568 = pi151 & ~pi191;
  assign n7569 = ~pi152 & pi192;
  assign n7570 = pi152 & ~pi192;
  assign n7571 = ~pi153 & pi193;
  assign n7572 = pi153 & ~pi193;
  assign n7573 = ~pi154 & pi194;
  assign n7574 = pi154 & ~pi194;
  assign n7575 = ~pi155 & pi195;
  assign n7576 = pi155 & ~pi195;
  assign n7577 = ~pi156 & pi196;
  assign n7578 = pi156 & ~pi196;
  assign n7579 = pi158 & ~pi198;
  assign n7580 = pi157 & ~pi197;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~pi157 & pi197;
  assign n7583 = ~n7581 & ~n7582;
  assign n7584 = ~n7578 & ~n7583;
  assign n7585 = ~n7577 & ~n7584;
  assign n7586 = ~n7576 & ~n7585;
  assign n7587 = ~n7575 & ~n7586;
  assign n7588 = ~n7574 & ~n7587;
  assign n7589 = ~n7573 & ~n7588;
  assign n7590 = ~n7572 & ~n7589;
  assign n7591 = ~n7571 & ~n7590;
  assign n7592 = ~n7570 & ~n7591;
  assign n7593 = ~n7569 & ~n7592;
  assign n7594 = ~n7568 & ~n7593;
  assign n7595 = ~n7567 & ~n7594;
  assign n7596 = ~n7566 & ~n7595;
  assign n7597 = n7537 & n7596;
  assign n7598 = ~n3283 & ~n3431;
  assign n7599 = ~n2721 & ~n2812;
  assign n7600 = n7598 & n7599;
  assign n7601 = n3819 & n4788;
  assign n7602 = n7600 & n7601;
  assign n7603 = n6181 & ~n6551;
  assign n7604 = ~n4281 & ~n5317;
  assign n7605 = n5732 & n7604;
  assign n7606 = n7603 & n7605;
  assign n7607 = n7602 & n7606;
  assign n7608 = n3808 & n7282;
  assign n7609 = ~n3285 & ~n3404;
  assign n7610 = n5722 & n7609;
  assign n7611 = ~n2664 & ~n2785;
  assign n7612 = n3810 & n7611;
  assign n7613 = n7610 & n7612;
  assign n7614 = ~n4254 & ~n5290;
  assign n7615 = ~n6144 & ~n6524;
  assign n7616 = n7614 & n7615;
  assign n7617 = n5721 & n7616;
  assign n7618 = n7613 & n7617;
  assign n7619 = pi015 & ~n501;
  assign n7620 = ~n504 & ~n1116;
  assign n7621 = n5713 & n7620;
  assign n7622 = n7619 & n7621;
  assign n7623 = ~n566 & ~n1374;
  assign n7624 = n5717 & n7623;
  assign n7625 = n3813 & n7624;
  assign n7626 = n7622 & n7625;
  assign n7627 = n7618 & n7626;
  assign n7628 = ~n1172 & n7627;
  assign n7629 = ~n1143 & n7628;
  assign n7630 = ~n996 & n7629;
  assign n7631 = ~n2306 & n7630;
  assign n7632 = ~n500 & n7631;
  assign n7633 = n2316 & n7632;
  assign n7634 = n7608 & n7633;
  assign n7635 = ~pi151 & pi271;
  assign n7636 = pi153 & ~pi273;
  assign n7637 = ~pi154 & pi274;
  assign n7638 = pi154 & ~pi274;
  assign n7639 = ~pi155 & pi275;
  assign n7640 = pi155 & ~pi275;
  assign n7641 = ~pi156 & pi276;
  assign n7642 = pi156 & ~pi276;
  assign n7643 = pi158 & ~pi278;
  assign n7644 = pi157 & ~pi277;
  assign n7645 = ~n7643 & ~n7644;
  assign n7646 = ~pi157 & pi277;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = ~n7642 & ~n7647;
  assign n7649 = ~n7641 & ~n7648;
  assign n7650 = ~n7640 & ~n7649;
  assign n7651 = ~n7639 & ~n7650;
  assign n7652 = ~n7638 & ~n7651;
  assign n7653 = ~n7637 & ~n7652;
  assign n7654 = ~n7636 & ~n7653;
  assign n7655 = ~pi153 & pi273;
  assign n7656 = ~pi152 & pi272;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = ~n7654 & n7657;
  assign n7659 = pi151 & ~pi271;
  assign n7660 = pi152 & ~pi272;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7658 & n7661;
  assign n7663 = ~n7635 & ~n7662;
  assign n7664 = ~pi151 & pi255;
  assign n7665 = pi153 & ~pi257;
  assign n7666 = ~pi154 & pi258;
  assign n7667 = pi154 & ~pi258;
  assign n7668 = ~pi155 & pi259;
  assign n7669 = pi155 & ~pi259;
  assign n7670 = ~pi156 & pi260;
  assign n7671 = pi156 & ~pi260;
  assign n7672 = pi158 & ~pi262;
  assign n7673 = pi157 & ~pi261;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = ~pi157 & pi261;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = ~n7671 & ~n7676;
  assign n7678 = ~n7670 & ~n7677;
  assign n7679 = ~n7669 & ~n7678;
  assign n7680 = ~n7668 & ~n7679;
  assign n7681 = ~n7667 & ~n7680;
  assign n7682 = ~n7666 & ~n7681;
  assign n7683 = ~n7665 & ~n7682;
  assign n7684 = ~pi153 & pi257;
  assign n7685 = ~pi152 & pi256;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = ~n7683 & n7686;
  assign n7688 = pi151 & ~pi255;
  assign n7689 = pi152 & ~pi256;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 = ~n7687 & n7690;
  assign n7692 = ~n7664 & ~n7691;
  assign n7693 = ~n7663 & ~n7692;
  assign n7694 = ~pi151 & pi231;
  assign n7695 = pi153 & ~pi233;
  assign n7696 = ~pi154 & pi234;
  assign n7697 = pi154 & ~pi234;
  assign n7698 = ~pi155 & pi235;
  assign n7699 = pi155 & ~pi235;
  assign n7700 = ~pi156 & pi236;
  assign n7701 = pi156 & ~pi236;
  assign n7702 = pi158 & ~pi238;
  assign n7703 = pi157 & ~pi237;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = ~pi157 & pi237;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = ~n7701 & ~n7706;
  assign n7708 = ~n7700 & ~n7707;
  assign n7709 = ~n7699 & ~n7708;
  assign n7710 = ~n7698 & ~n7709;
  assign n7711 = ~n7697 & ~n7710;
  assign n7712 = ~n7696 & ~n7711;
  assign n7713 = ~n7695 & ~n7712;
  assign n7714 = ~pi153 & pi233;
  assign n7715 = ~pi152 & pi232;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = ~n7713 & n7716;
  assign n7718 = pi151 & ~pi231;
  assign n7719 = pi152 & ~pi232;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = ~n7717 & n7720;
  assign n7722 = ~n7694 & ~n7721;
  assign n7723 = ~pi151 & pi239;
  assign n7724 = pi153 & ~pi241;
  assign n7725 = ~pi154 & pi242;
  assign n7726 = pi154 & ~pi242;
  assign n7727 = ~pi155 & pi243;
  assign n7728 = pi155 & ~pi243;
  assign n7729 = ~pi156 & pi244;
  assign n7730 = pi156 & ~pi244;
  assign n7731 = pi158 & ~pi246;
  assign n7732 = pi157 & ~pi245;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = ~pi157 & pi245;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = ~n7730 & ~n7735;
  assign n7737 = ~n7729 & ~n7736;
  assign n7738 = ~n7728 & ~n7737;
  assign n7739 = ~n7727 & ~n7738;
  assign n7740 = ~n7726 & ~n7739;
  assign n7741 = ~n7725 & ~n7740;
  assign n7742 = ~n7724 & ~n7741;
  assign n7743 = ~pi153 & pi241;
  assign n7744 = ~pi152 & pi240;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = ~n7742 & n7745;
  assign n7747 = pi151 & ~pi239;
  assign n7748 = pi152 & ~pi240;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = ~n7746 & n7749;
  assign n7751 = ~n7723 & ~n7750;
  assign n7752 = ~n7722 & ~n7751;
  assign n7753 = n7693 & n7752;
  assign n7754 = ~n7240 & ~n7277;
  assign n7755 = ~n1402 & ~n7754;
  assign n7756 = n4786 & n7755;
  assign n7757 = n7753 & n7756;
  assign n7758 = n7634 & n7757;
  assign n7759 = n7607 & n7758;
  assign n7760 = n7597 & n7759;
  assign n7761 = ~n6137 & n7760;
  assign n7762 = n6193 & n7761;
  assign n7763 = n6134 & n7762;
  assign n7764 = ~n7298 & ~n7763;
  assign n7765 = ~n7211 & n7764;
  assign po008 = n7205 | ~n7765;
  assign n7767 = n6872 & ~n7073;
  assign n7768 = n3089 & n5835;
  assign n7769 = n1680 & n3085;
  assign n7770 = n3883 & n7769;
  assign n7771 = n5810 & n7770;
  assign n7772 = n7768 & n7771;
  assign n7773 = ~n6838 & n7772;
  assign n7774 = ~n2242 & n7773;
  assign n7775 = ~n3095 & n7774;
  assign n7776 = ~n3997 & n7775;
  assign n7777 = ~n4003 & n7776;
  assign n7778 = ~n4837 & n7777;
  assign n7779 = ~n5822 & n7778;
  assign n7780 = ~n6837 & n7779;
  assign n7781 = ~n6820 & n7780;
  assign n7782 = ~n6836 & n7781;
  assign n7783 = n6857 & n7782;
  assign n7784 = n6835 & n7783;
  assign n7785 = n6830 & n7784;
  assign n7786 = n6864 & ~n7785;
  assign n7787 = ~n7767 & ~n7786;
  assign n7788 = n6869 & ~n7204;
  assign n7789 = ~n1026 & n6723;
  assign n7790 = n6787 & n7789;
  assign n7791 = n1239 & n7790;
  assign n7792 = ~n1270 & n7791;
  assign n7793 = n844 & n7792;
  assign n7794 = ~n1372 & n7793;
  assign n7795 = ~n2243 & n7794;
  assign n7796 = ~n6785 & n7795;
  assign n7797 = ~n3104 & n7796;
  assign n7798 = ~n3971 & n7797;
  assign n7799 = ~n4003 & n7798;
  assign n7800 = ~n4872 & n7799;
  assign n7801 = ~n5801 & n7800;
  assign n7802 = ~n6761 & n7801;
  assign n7803 = ~n6760 & n7802;
  assign n7804 = ~n6759 & n7803;
  assign n7805 = n6822 & n7804;
  assign n7806 = n6758 & n7805;
  assign n7807 = n6722 & n7806;
  assign n7808 = n6889 & ~n7807;
  assign n7809 = ~n7788 & ~n7808;
  assign n7810 = n7787 & n7809;
  assign n7811 = n4847 & n5718;
  assign n7812 = n3941 & n5722;
  assign n7813 = n3859 & n5754;
  assign n7814 = n7812 & n7813;
  assign n7815 = n6740 & ~n7240;
  assign n7816 = n4849 & n5757;
  assign n7817 = n7815 & n7816;
  assign n7818 = n7814 & n7817;
  assign n7819 = n7811 & n7818;
  assign n7820 = ~n1172 & n7819;
  assign n7821 = ~n996 & n7820;
  assign n7822 = ~n2306 & n7821;
  assign n7823 = ~n500 & n7822;
  assign n7824 = n6677 & n7823;
  assign n7825 = n7280 & n7824;
  assign n7826 = n7284 & n7825;
  assign n7827 = ~n7236 & n7826;
  assign n7828 = ~n6137 & n7827;
  assign n7829 = n6193 & n7828;
  assign n7830 = n6134 & n7829;
  assign n7831 = ~n7235 & n7830;
  assign n7832 = n7296 & n7831;
  assign po161 = n7231 & n7832;
  assign n7834 = n3053 & ~po161;
  assign n7835 = n6867 & ~n7029;
  assign n7836 = ~n7834 & ~n7835;
  assign n7837 = n6868 & ~n6967;
  assign n7838 = n6888 & ~n7095;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7836 & n7839;
  assign n7841 = n6862 & ~n6951;
  assign n7842 = n6873 & ~n6917;
  assign n7843 = ~n3256 & ~n3404;
  assign n7844 = n6762 & n7843;
  assign n7845 = n3941 & n7611;
  assign n7846 = n7844 & n7845;
  assign n7847 = ~n6524 & n6740;
  assign n7848 = n5757 & n7614;
  assign n7849 = n7847 & n7848;
  assign n7850 = n7846 & n7849;
  assign n7851 = n2246 & n7621;
  assign n7852 = ~n1374 & ~n1435;
  assign n7853 = n3859 & n7852;
  assign n7854 = n5718 & n7853;
  assign n7855 = n7851 & n7854;
  assign n7856 = n7850 & n7855;
  assign n7857 = ~n1172 & n7856;
  assign n7858 = ~n1143 & n7857;
  assign n7859 = ~n996 & n7858;
  assign n7860 = ~n2306 & n7859;
  assign n7861 = ~n500 & n7860;
  assign n7862 = n2316 & n7861;
  assign n7863 = n7608 & n7862;
  assign n7864 = n7757 & n7863;
  assign n7865 = n7607 & n7864;
  assign n7866 = n7597 & n7865;
  assign n7867 = ~n6137 & n7866;
  assign n7868 = n6193 & n7867;
  assign n7869 = n6134 & n7868;
  assign n7870 = n2813 & ~n7869;
  assign n7871 = n2784 & n3838;
  assign n7872 = ~n3024 & n7871;
  assign n7873 = ~n2934 & n7872;
  assign n7874 = n2634 & n7873;
  assign n7875 = ~n3066 & n7874;
  assign n7876 = ~n3983 & n7875;
  assign n7877 = ~n4003 & n7876;
  assign n7878 = ~n4024 & n7877;
  assign n7879 = ~n4999 & n7878;
  assign n7880 = ~n5827 & n7879;
  assign n7881 = ~n7870 & n7880;
  assign n7882 = ~n7842 & n7881;
  assign n7883 = ~n6893 & n7882;
  assign n7884 = ~n7841 & n7883;
  assign n7885 = n6863 & ~n7014;
  assign n7886 = n6874 & ~n7158;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = n7884 & n7887;
  assign n7889 = n7840 & n7888;
  assign n7890 = n7810 & n7889;
  assign n7891 = n6855 & ~n7073;
  assign n7892 = n6827 & ~n6893;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = n6833 & ~n7204;
  assign n7895 = n6826 & ~n7807;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = n7893 & n7896;
  assign n7898 = n1804 & ~po161;
  assign n7899 = n6831 & ~n7029;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = n6832 & ~n6967;
  assign n7902 = n6856 & ~n7095;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = n7900 & n7903;
  assign n7905 = n6836 & ~n6951;
  assign n7906 = n6837 & ~n6917;
  assign n7907 = n1403 & ~n7869;
  assign n7908 = ~n1958 & n3889;
  assign n7909 = ~n1617 & n3069;
  assign n7910 = n6842 & n7909;
  assign n7911 = n7908 & n7910;
  assign n7912 = ~n2242 & n7911;
  assign n7913 = ~n3095 & n7912;
  assign n7914 = ~n3997 & n7913;
  assign n7915 = ~n4003 & n7914;
  assign n7916 = ~n4837 & n7915;
  assign n7917 = ~n5822 & n7916;
  assign n7918 = ~n6820 & n7917;
  assign n7919 = ~n7907 & n7918;
  assign n7920 = ~n7906 & n7919;
  assign n7921 = ~n7785 & n7920;
  assign n7922 = ~n7905 & n7921;
  assign n7923 = n6828 & ~n7014;
  assign n7924 = n6838 & ~n7158;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = n7922 & n7925;
  assign n7927 = n7904 & n7926;
  assign n7928 = n7897 & n7927;
  assign n7929 = n6719 & ~n7014;
  assign n7930 = n6785 & ~n7158;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = n6759 & ~n7073;
  assign n7933 = n6821 & ~n7785;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = n7931 & n7934;
  assign n7936 = n1299 & ~po161;
  assign n7937 = n6756 & ~n7029;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = n6760 & ~n6967;
  assign n7940 = n6803 & ~n7095;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = n7938 & n7941;
  assign n7943 = n6720 & ~n6893;
  assign n7944 = n6761 & ~n6917;
  assign n7945 = n1144 & ~n7869;
  assign n7946 = pi001 & ~n1115;
  assign n7947 = ~n1026 & n7946;
  assign n7948 = ~n1086 & n7947;
  assign n7949 = n1239 & n7948;
  assign n7950 = ~n1270 & n7949;
  assign n7951 = n844 & n7950;
  assign n7952 = ~n1372 & n7951;
  assign n7953 = ~n2243 & n7952;
  assign n7954 = ~n3104 & n7953;
  assign n7955 = ~n3971 & n7954;
  assign n7956 = ~n4003 & n7955;
  assign n7957 = ~n4872 & n7956;
  assign n7958 = ~n5801 & n7957;
  assign n7959 = ~n6739 & n7958;
  assign n7960 = ~n7945 & n7959;
  assign n7961 = ~n7944 & n7960;
  assign n7962 = ~n7807 & n7961;
  assign n7963 = ~n7943 & n7962;
  assign n7964 = n6755 & ~n7204;
  assign n7965 = n6718 & ~n6951;
  assign n7966 = ~n7964 & ~n7965;
  assign n7967 = n7963 & n7966;
  assign n7968 = n7942 & n7967;
  assign n7969 = n7935 & n7968;
  assign n7970 = ~n7928 & ~n7969;
  assign n7971 = ~n7890 & n7970;
  assign n7972 = ~pi005 & ~n2543;
  assign n7973 = n5772 & n7972;
  assign n7974 = ~n2783 & ~n2842;
  assign n7975 = ~n2663 & n7974;
  assign n7976 = n5775 & n7975;
  assign n7977 = ~n2934 & ~n3024;
  assign n7978 = n7976 & n7977;
  assign n7979 = n7973 & n7978;
  assign n7980 = ~n3066 & n7979;
  assign n7981 = ~n3983 & n7980;
  assign n7982 = ~n4003 & n7981;
  assign n7983 = ~n4024 & n7982;
  assign n7984 = ~n4999 & n7983;
  assign n7985 = ~n5827 & n7984;
  assign n7986 = ~n7870 & n7985;
  assign n7987 = ~n7842 & n7986;
  assign n7988 = ~n6893 & n7987;
  assign n7989 = ~n7841 & n7988;
  assign n7990 = n7887 & n7989;
  assign n7991 = n7840 & n7990;
  assign n7992 = n7810 & n7991;
  assign n7993 = n6911 & ~n7785;
  assign n7994 = n6912 & ~n6917;
  assign n7995 = ~n7993 & n7994;
  assign n7996 = n6915 & ~n7807;
  assign n7997 = ~n6893 & n6914;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = n7995 & n7998;
  assign n8000 = ~n7992 & ~n7999;
  assign n8001 = ~n7971 & n8000;
  assign n8002 = n6932 & ~n7158;
  assign n8003 = ~n6893 & n6920;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = n6921 & ~n7785;
  assign n8006 = n6922 & ~n7807;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = n8004 & n8007;
  assign n8009 = n3136 & ~po161;
  assign n8010 = n6926 & ~n7029;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = n6925 & ~n6967;
  assign n8013 = n6947 & ~n7095;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = n8011 & n8014;
  assign n8016 = n6930 & ~n7014;
  assign n8017 = ~n6917 & n6931;
  assign n8018 = n3432 & ~n7869;
  assign n8019 = n4096 & n6935;
  assign n8020 = n4104 & n8019;
  assign n8021 = ~n3464 & n4101;
  assign n8022 = ~n3165 & n8021;
  assign n8023 = n8020 & n8022;
  assign n8024 = ~n3940 & n8023;
  assign n8025 = ~n4001 & n8024;
  assign n8026 = ~n5043 & n8025;
  assign n8027 = ~n5943 & n8026;
  assign n8028 = ~n8018 & n8027;
  assign n8029 = ~n8017 & n8028;
  assign n8030 = ~n6951 & n8029;
  assign n8031 = ~n8016 & n8030;
  assign n8032 = n6927 & ~n7204;
  assign n8033 = n6946 & ~n7073;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 = n8031 & n8034;
  assign n8036 = n8015 & n8035;
  assign n8037 = n8008 & n8036;
  assign n8038 = ~n5917 & n5969;
  assign n8039 = ~n6917 & n8038;
  assign n8040 = ~n7993 & n8039;
  assign n8041 = n7998 & n8040;
  assign n8042 = ~n8037 & ~n8041;
  assign n8043 = ~n8001 & n8042;
  assign n8044 = ~n6893 & n6962;
  assign n8045 = n6959 & ~n6967;
  assign n8046 = ~n8017 & n8045;
  assign n8047 = ~n8044 & n8046;
  assign n8048 = n6963 & ~n7785;
  assign n8049 = ~n6951 & n6958;
  assign n8050 = n6964 & ~n7807;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = ~n8048 & n8051;
  assign n8053 = n8047 & n8052;
  assign n8054 = ~pi007 & ~n3524;
  assign n8055 = n3800 & n8054;
  assign n8056 = n3374 & ~n3403;
  assign n8057 = n3681 & n8056;
  assign n8058 = ~n3165 & ~n3464;
  assign n8059 = n8057 & n8058;
  assign n8060 = n8055 & n8059;
  assign n8061 = ~n3940 & n8060;
  assign n8062 = ~n4001 & n8061;
  assign n8063 = ~n5043 & n8062;
  assign n8064 = ~n5943 & n8063;
  assign n8065 = ~n8018 & n8064;
  assign n8066 = ~n8017 & n8065;
  assign n8067 = ~n6951 & n8066;
  assign n8068 = ~n8016 & n8067;
  assign n8069 = n8034 & n8068;
  assign n8070 = n8015 & n8069;
  assign n8071 = n8008 & n8070;
  assign n8072 = ~n8053 & ~n8071;
  assign n8073 = ~n8043 & n8072;
  assign n8074 = ~n5058 & n5077;
  assign n8075 = ~n5967 & n8074;
  assign n8076 = ~n6967 & n8075;
  assign n8077 = ~n8017 & n8076;
  assign n8078 = ~n8044 & n8077;
  assign n8079 = n8052 & n8078;
  assign n8080 = ~n6951 & n6987;
  assign n8081 = ~n6893 & n7010;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = n6996 & ~n7785;
  assign n8084 = n7009 & ~n7807;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = n8082 & n8085;
  assign n8087 = n6988 & ~n7095;
  assign n8088 = ~n8045 & ~n8087;
  assign n8089 = n6992 & ~n7029;
  assign n8090 = n4521 & ~po161;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = n8088 & n8091;
  assign n8093 = n6989 & ~n7073;
  assign n8094 = n4282 & ~n7869;
  assign n8095 = ~n4311 & ~n4489;
  assign n8096 = n5084 & n8095;
  assign n8097 = n5083 & n5087;
  assign n8098 = n8096 & n8097;
  assign n8099 = ~n4163 & n7032;
  assign n8100 = ~n4192 & n8099;
  assign n8101 = n8098 & n8100;
  assign n8102 = ~n4817 & n8101;
  assign n8103 = ~n4902 & n8102;
  assign n8104 = ~n6001 & n8103;
  assign n8105 = ~n8094 & n8104;
  assign n8106 = ~n8017 & n8105;
  assign n8107 = ~n7014 & n8106;
  assign n8108 = ~n8093 & n8107;
  assign n8109 = n6993 & ~n7204;
  assign n8110 = n6997 & ~n7158;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = n8108 & n8111;
  assign n8113 = n8092 & n8112;
  assign n8114 = n8086 & n8113;
  assign n8115 = ~n8079 & ~n8114;
  assign n8116 = ~n8073 & n8115;
  assign n8117 = ~pi009 & ~n4677;
  assign n8118 = n7030 & n8117;
  assign n8119 = n4490 & n5094;
  assign n8120 = n6999 & n8119;
  assign n8121 = n4193 & n8120;
  assign n8122 = n8118 & n8121;
  assign n8123 = ~n4817 & n8122;
  assign n8124 = ~n4902 & n8123;
  assign n8125 = ~n6001 & n8124;
  assign n8126 = ~n8094 & n8125;
  assign n8127 = ~n8017 & n8126;
  assign n8128 = ~n7014 & n8127;
  assign n8129 = ~n8093 & n8128;
  assign n8130 = n8111 & n8129;
  assign n8131 = n8092 & n8130;
  assign n8132 = n8086 & n8131;
  assign n8133 = ~n6893 & n7025;
  assign n8134 = ~n6951 & n7019;
  assign n8135 = n7026 & ~n7807;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = ~n8133 & n8136;
  assign n8138 = n7022 & ~n7029;
  assign n8139 = ~n8017 & n8138;
  assign n8140 = ~n8045 & n8139;
  assign n8141 = ~n7014 & n7017;
  assign n8142 = n7018 & ~n7785;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = n8140 & n8143;
  assign n8145 = n8137 & n8144;
  assign n8146 = ~n8132 & ~n8145;
  assign n8147 = ~n8116 & n8146;
  assign n8148 = n7057 & ~n7158;
  assign n8149 = ~n6893 & n7056;
  assign n8150 = ~n8148 & ~n8149;
  assign n8151 = n7069 & ~n7807;
  assign n8152 = n7050 & ~n7785;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n8150 & n8153;
  assign n8155 = ~n8045 & ~n8138;
  assign n8156 = n5199 & ~po161;
  assign n8157 = n7049 & ~n7095;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = n8155 & n8158;
  assign n8160 = ~n7014 & n7068;
  assign n8161 = n5318 & ~n7869;
  assign n8162 = n5439 & n5688;
  assign n8163 = ~n5289 & ~n5527;
  assign n8164 = n5260 & n8163;
  assign n8165 = ~n5469 & n8164;
  assign n8166 = ~n5170 & n8165;
  assign n8167 = n8162 & n8166;
  assign n8168 = ~n5808 & n8167;
  assign n8169 = ~n6056 & n8168;
  assign n8170 = ~n8161 & n8169;
  assign n8171 = ~n8017 & n8170;
  assign n8172 = ~n7073 & n8171;
  assign n8173 = ~n8160 & n8172;
  assign n8174 = n7053 & ~n7204;
  assign n8175 = ~n6951 & n7048;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = n8173 & n8176;
  assign n8178 = n8159 & n8177;
  assign n8179 = n8154 & n8178;
  assign n8180 = ~n4881 & n5107;
  assign n8181 = ~n6027 & n8180;
  assign n8182 = ~n7029 & n8181;
  assign n8183 = ~n8017 & n8182;
  assign n8184 = ~n8045 & n8183;
  assign n8185 = n8143 & n8184;
  assign n8186 = n8137 & n8185;
  assign n8187 = ~n8179 & ~n8186;
  assign n8188 = ~n8147 & n8187;
  assign n8189 = ~pi011 & ~n5598;
  assign n8190 = n7096 & n8189;
  assign n8191 = ~n5527 & n6074;
  assign n8192 = n7099 & n8191;
  assign n8193 = n6036 & n8192;
  assign n8194 = n8190 & n8193;
  assign n8195 = ~n5808 & n8194;
  assign n8196 = ~n6056 & n8195;
  assign n8197 = ~n8161 & n8196;
  assign n8198 = ~n8017 & n8197;
  assign n8199 = ~n7073 & n8198;
  assign n8200 = ~n8160 & n8199;
  assign n8201 = n8176 & n8200;
  assign n8202 = n8159 & n8201;
  assign n8203 = n8154 & n8202;
  assign n8204 = ~n6951 & n7082;
  assign n8205 = ~n7073 & n7081;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = ~n6893 & n7085;
  assign n8208 = n7092 & ~n7807;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = n8206 & n8209;
  assign n8211 = ~n7095 & n7152;
  assign n8212 = ~n8017 & n8211;
  assign n8213 = n8155 & n8212;
  assign n8214 = n7091 & ~n7785;
  assign n8215 = ~n7014 & n7084;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = n8213 & n8216;
  assign n8218 = n8210 & n8217;
  assign n8219 = ~n8203 & ~n8218;
  assign n8220 = ~n8188 & n8219;
  assign n8221 = ~n6893 & n7130;
  assign n8222 = ~n7073 & n7154;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = n7141 & ~n7204;
  assign n8225 = n7118 & ~n7785;
  assign n8226 = ~n8224 & ~n8225;
  assign n8227 = n8223 & n8226;
  assign n8228 = n6253 & ~po161;
  assign n8229 = ~n8211 & ~n8228;
  assign n8230 = n8155 & n8229;
  assign n8231 = ~n6951 & n7150;
  assign n8232 = n6552 & ~n7869;
  assign n8233 = n6402 & n6614;
  assign n8234 = n6343 & n6462;
  assign n8235 = n8233 & n8234;
  assign n8236 = n6523 & n6673;
  assign n8237 = ~n6282 & n8236;
  assign n8238 = ~n6224 & n8237;
  assign n8239 = n8235 & n8238;
  assign n8240 = ~n6784 & n8239;
  assign n8241 = ~n8232 & n8240;
  assign n8242 = ~n8017 & n8241;
  assign n8243 = ~n7158 & n8242;
  assign n8244 = ~n8231 & n8243;
  assign n8245 = ~n7014 & n7146;
  assign n8246 = n7125 & ~n7807;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n8244 & n8247;
  assign n8249 = n8230 & n8248;
  assign n8250 = n8227 & n8249;
  assign n8251 = ~n6114 & n6116;
  assign n8252 = ~n7095 & n8251;
  assign n8253 = ~n8017 & n8252;
  assign n8254 = n8155 & n8253;
  assign n8255 = n8216 & n8254;
  assign n8256 = n8210 & n8255;
  assign n8257 = ~n8250 & ~n8256;
  assign n8258 = ~n8220 & n8257;
  assign n8259 = ~pi013 & ~n6432;
  assign n8260 = n7170 & n8259;
  assign n8261 = ~n6522 & n7172;
  assign n8262 = n7177 & n8261;
  assign n8263 = ~n6224 & ~n6282;
  assign n8264 = n8262 & n8263;
  assign n8265 = n8260 & n8264;
  assign n8266 = ~n6784 & n8265;
  assign n8267 = ~n8232 & n8266;
  assign n8268 = ~n8017 & n8267;
  assign n8269 = ~n7158 & n8268;
  assign n8270 = ~n8231 & n8269;
  assign n8271 = n8247 & n8270;
  assign n8272 = n8230 & n8271;
  assign n8273 = n8227 & n8272;
  assign n8274 = ~n6893 & n7197;
  assign n8275 = ~n7014 & n7199;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n7158 & n7193;
  assign n8278 = ~n7073 & n7190;
  assign n8279 = ~n8277 & ~n8278;
  assign n8280 = n8276 & n8279;
  assign n8281 = n8155 & ~n8211;
  assign n8282 = ~n6951 & n7188;
  assign n8283 = ~n6754 & ~n8017;
  assign n8284 = ~n7204 & n8283;
  assign n8285 = ~n8282 & n8284;
  assign n8286 = n7200 & ~n7807;
  assign n8287 = n7189 & ~n7785;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = n8285 & n8288;
  assign n8290 = n8281 & n8289;
  assign n8291 = n8280 & n8290;
  assign n8292 = ~n2813 & ~n3066;
  assign n8293 = ~n3983 & n8292;
  assign n8294 = ~n4024 & n8293;
  assign n8295 = ~n4999 & n8294;
  assign n8296 = ~n5827 & n8295;
  assign n8297 = ~n6893 & n8296;
  assign n8298 = ~n6552 & ~n6784;
  assign n8299 = ~n7158 & n8298;
  assign n8300 = ~n3432 & ~n3940;
  assign n8301 = ~n4001 & n8300;
  assign n8302 = ~n5043 & n8301;
  assign n8303 = ~n5943 & n8302;
  assign n8304 = ~n6951 & n8303;
  assign n8305 = ~n8299 & ~n8304;
  assign n8306 = ~n8297 & n8305;
  assign n8307 = ~n1403 & ~n2242;
  assign n8308 = ~n3095 & n8307;
  assign n8309 = ~n3997 & n8308;
  assign n8310 = ~n4837 & n8309;
  assign n8311 = ~n5822 & n8310;
  assign n8312 = ~n6820 & n8311;
  assign n8313 = ~n7785 & n8312;
  assign n8314 = ~n6754 & ~n7204;
  assign n8315 = ~n8313 & ~n8314;
  assign n8316 = ~n1144 & ~n1372;
  assign n8317 = ~n2243 & n8316;
  assign n8318 = ~n3104 & n8317;
  assign n8319 = ~n3971 & n8318;
  assign n8320 = ~n4872 & n8319;
  assign n8321 = ~n5801 & n8320;
  assign n8322 = ~n6739 & n8321;
  assign n8323 = ~n7807 & n8322;
  assign n8324 = ~n5318 & ~n5808;
  assign n8325 = ~n6056 & n8324;
  assign n8326 = ~n7073 & n8325;
  assign n8327 = ~n8323 & ~n8326;
  assign n8328 = n8315 & n8327;
  assign n8329 = n7754 & ~po161;
  assign n8330 = ~n8138 & ~n8211;
  assign n8331 = ~n8329 & n8330;
  assign n8332 = ~n4282 & ~n4817;
  assign n8333 = ~n4902 & n8332;
  assign n8334 = ~n6001 & n8333;
  assign n8335 = ~n7014 & n8334;
  assign n8336 = n7536 & n7753;
  assign n8337 = n7417 & ~n7566;
  assign n8338 = ~n7595 & n8337;
  assign n8339 = n8336 & n8338;
  assign n8340 = ~n7869 & n8339;
  assign n8341 = ~n8017 & n8340;
  assign n8342 = ~n8045 & n8341;
  assign n8343 = ~n8335 & n8342;
  assign n8344 = n8331 & n8343;
  assign n8345 = n8328 & n8344;
  assign n8346 = n8306 & n8345;
  assign n8347 = ~n8291 & ~n8346;
  assign n8348 = ~n8273 & n8347;
  assign n8349 = ~n8258 & n8348;
  assign n8350 = pi014 & ~n6754;
  assign n8351 = ~n8017 & n8350;
  assign n8352 = ~n7204 & n8351;
  assign n8353 = ~n8282 & n8352;
  assign n8354 = n8288 & n8353;
  assign n8355 = n8281 & n8354;
  assign n8356 = n8280 & n8355;
  assign n8357 = pi015 & ~n7663;
  assign n8358 = ~n7692 & ~n7722;
  assign n8359 = ~n7446 & ~n7751;
  assign n8360 = n8358 & n8359;
  assign n8361 = n8357 & n8360;
  assign n8362 = ~n7356 & ~n7386;
  assign n8363 = ~n7415 & n8362;
  assign n8364 = ~n7475 & ~n7505;
  assign n8365 = ~n7327 & ~n7534;
  assign n8366 = n8364 & n8365;
  assign n8367 = n8363 & n8366;
  assign n8368 = n7596 & n8367;
  assign n8369 = n8361 & n8368;
  assign n8370 = ~n7869 & n8369;
  assign n8371 = ~n8017 & n8370;
  assign n8372 = ~n8045 & n8371;
  assign n8373 = ~n8335 & n8372;
  assign n8374 = n8331 & n8373;
  assign n8375 = n8328 & n8374;
  assign n8376 = n8306 & n8375;
  assign n8377 = ~n8356 & ~n8376;
  assign n8378 = ~n8349 & n8377;
  assign n8379 = ~n7158 & n7236;
  assign n8380 = ~n7014 & n7293;
  assign n8381 = ~n6951 & n7235;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = ~n8379 & n8382;
  assign n8384 = ~n7073 & n7295;
  assign n8385 = ~n6893 & n7223;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n7229 & ~n7785;
  assign n8388 = n7218 & ~n7807;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = n8386 & n8389;
  assign n8391 = ~n7754 & ~n7869;
  assign n8392 = ~po161 & ~n8391;
  assign n8393 = ~n8017 & n8392;
  assign n8394 = ~n8314 & n8393;
  assign n8395 = n8281 & n8394;
  assign n8396 = n8390 & n8395;
  assign n8397 = n8383 & n8396;
  assign n8398 = ~pi167 & pi191;
  assign n8399 = pi167 & ~pi191;
  assign n8400 = ~pi168 & pi192;
  assign n8401 = pi168 & ~pi192;
  assign n8402 = ~pi169 & pi193;
  assign n8403 = pi169 & ~pi193;
  assign n8404 = ~pi170 & pi194;
  assign n8405 = pi170 & ~pi194;
  assign n8406 = ~pi171 & pi195;
  assign n8407 = pi171 & ~pi195;
  assign n8408 = ~pi172 & pi196;
  assign n8409 = pi172 & ~pi196;
  assign n8410 = pi174 & ~pi198;
  assign n8411 = pi173 & ~pi197;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = ~pi173 & pi197;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = ~n8409 & ~n8414;
  assign n8416 = ~n8408 & ~n8415;
  assign n8417 = ~n8407 & ~n8416;
  assign n8418 = ~n8406 & ~n8417;
  assign n8419 = ~n8405 & ~n8418;
  assign n8420 = ~n8404 & ~n8419;
  assign n8421 = ~n8403 & ~n8420;
  assign n8422 = ~n8402 & ~n8421;
  assign n8423 = ~n8401 & ~n8422;
  assign n8424 = ~n8400 & ~n8423;
  assign n8425 = ~n8399 & ~n8424;
  assign n8426 = ~n8398 & ~n8425;
  assign n8427 = ~pi167 & pi263;
  assign n8428 = pi169 & ~pi265;
  assign n8429 = ~pi170 & pi266;
  assign n8430 = pi170 & ~pi266;
  assign n8431 = ~pi171 & pi267;
  assign n8432 = pi171 & ~pi267;
  assign n8433 = ~pi172 & pi268;
  assign n8434 = pi172 & ~pi268;
  assign n8435 = pi174 & ~pi270;
  assign n8436 = pi173 & ~pi269;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = ~pi173 & pi269;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = ~n8434 & ~n8439;
  assign n8441 = ~n8433 & ~n8440;
  assign n8442 = ~n8432 & ~n8441;
  assign n8443 = ~n8431 & ~n8442;
  assign n8444 = ~n8430 & ~n8443;
  assign n8445 = ~n8429 & ~n8444;
  assign n8446 = ~n8428 & ~n8445;
  assign n8447 = ~pi169 & pi265;
  assign n8448 = ~pi168 & pi264;
  assign n8449 = ~n8447 & ~n8448;
  assign n8450 = ~n8446 & n8449;
  assign n8451 = pi167 & ~pi263;
  assign n8452 = pi168 & ~pi264;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = ~n8450 & n8453;
  assign n8455 = ~n8427 & ~n8454;
  assign n8456 = ~pi167 & pi255;
  assign n8457 = pi169 & ~pi257;
  assign n8458 = ~pi170 & pi258;
  assign n8459 = pi170 & ~pi258;
  assign n8460 = ~pi171 & pi259;
  assign n8461 = pi171 & ~pi259;
  assign n8462 = ~pi172 & pi260;
  assign n8463 = pi172 & ~pi260;
  assign n8464 = pi174 & ~pi262;
  assign n8465 = pi173 & ~pi261;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = ~pi173 & pi261;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = ~n8463 & ~n8468;
  assign n8470 = ~n8462 & ~n8469;
  assign n8471 = ~n8461 & ~n8470;
  assign n8472 = ~n8460 & ~n8471;
  assign n8473 = ~n8459 & ~n8472;
  assign n8474 = ~n8458 & ~n8473;
  assign n8475 = ~n8457 & ~n8474;
  assign n8476 = ~pi169 & pi257;
  assign n8477 = ~pi168 & pi256;
  assign n8478 = ~n8476 & ~n8477;
  assign n8479 = ~n8475 & n8478;
  assign n8480 = pi167 & ~pi255;
  assign n8481 = pi168 & ~pi256;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = ~n8479 & n8482;
  assign n8484 = ~n8456 & ~n8483;
  assign n8485 = ~n8455 & ~n8484;
  assign n8486 = ~pi167 & pi231;
  assign n8487 = pi169 & ~pi233;
  assign n8488 = ~pi170 & pi234;
  assign n8489 = pi170 & ~pi234;
  assign n8490 = ~pi171 & pi235;
  assign n8491 = pi171 & ~pi235;
  assign n8492 = ~pi172 & pi236;
  assign n8493 = pi172 & ~pi236;
  assign n8494 = pi174 & ~pi238;
  assign n8495 = pi173 & ~pi237;
  assign n8496 = ~n8494 & ~n8495;
  assign n8497 = ~pi173 & pi237;
  assign n8498 = ~n8496 & ~n8497;
  assign n8499 = ~n8493 & ~n8498;
  assign n8500 = ~n8492 & ~n8499;
  assign n8501 = ~n8491 & ~n8500;
  assign n8502 = ~n8490 & ~n8501;
  assign n8503 = ~n8489 & ~n8502;
  assign n8504 = ~n8488 & ~n8503;
  assign n8505 = ~n8487 & ~n8504;
  assign n8506 = ~pi169 & pi233;
  assign n8507 = ~pi168 & pi232;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = ~n8505 & n8508;
  assign n8510 = pi167 & ~pi231;
  assign n8511 = pi168 & ~pi232;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 = ~n8509 & n8512;
  assign n8514 = ~n8486 & ~n8513;
  assign n8515 = ~pi167 & pi239;
  assign n8516 = pi169 & ~pi241;
  assign n8517 = ~pi170 & pi242;
  assign n8518 = pi170 & ~pi242;
  assign n8519 = ~pi171 & pi243;
  assign n8520 = pi171 & ~pi243;
  assign n8521 = ~pi172 & pi244;
  assign n8522 = pi172 & ~pi244;
  assign n8523 = pi174 & ~pi246;
  assign n8524 = pi173 & ~pi245;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = ~pi173 & pi245;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~n8522 & ~n8527;
  assign n8529 = ~n8521 & ~n8528;
  assign n8530 = ~n8520 & ~n8529;
  assign n8531 = ~n8519 & ~n8530;
  assign n8532 = ~n8518 & ~n8531;
  assign n8533 = ~n8517 & ~n8532;
  assign n8534 = ~n8516 & ~n8533;
  assign n8535 = ~pi169 & pi241;
  assign n8536 = ~pi168 & pi240;
  assign n8537 = ~n8535 & ~n8536;
  assign n8538 = ~n8534 & n8537;
  assign n8539 = pi167 & ~pi239;
  assign n8540 = pi168 & ~pi240;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = ~n8538 & n8541;
  assign n8543 = ~n8515 & ~n8542;
  assign n8544 = ~n8514 & ~n8543;
  assign n8545 = n8485 & n8544;
  assign n8546 = ~pi167 & pi247;
  assign n8547 = pi169 & ~pi249;
  assign n8548 = ~pi170 & pi250;
  assign n8549 = pi170 & ~pi250;
  assign n8550 = ~pi171 & pi251;
  assign n8551 = pi171 & ~pi251;
  assign n8552 = ~pi172 & pi252;
  assign n8553 = pi172 & ~pi252;
  assign n8554 = pi174 & ~pi254;
  assign n8555 = pi173 & ~pi253;
  assign n8556 = ~n8554 & ~n8555;
  assign n8557 = ~pi173 & pi253;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = ~n8553 & ~n8558;
  assign n8560 = ~n8552 & ~n8559;
  assign n8561 = ~n8551 & ~n8560;
  assign n8562 = ~n8550 & ~n8561;
  assign n8563 = ~n8549 & ~n8562;
  assign n8564 = ~n8548 & ~n8563;
  assign n8565 = ~n8547 & ~n8564;
  assign n8566 = ~pi169 & pi249;
  assign n8567 = ~pi168 & pi248;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = ~n8565 & n8568;
  assign n8570 = pi167 & ~pi247;
  assign n8571 = pi168 & ~pi248;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = ~n8569 & n8572;
  assign n8574 = ~n8546 & ~n8573;
  assign n8575 = ~pi167 & pi215;
  assign n8576 = pi169 & ~pi217;
  assign n8577 = ~pi170 & pi218;
  assign n8578 = pi170 & ~pi218;
  assign n8579 = ~pi171 & pi219;
  assign n8580 = pi171 & ~pi219;
  assign n8581 = ~pi172 & pi220;
  assign n8582 = pi172 & ~pi220;
  assign n8583 = pi174 & ~pi222;
  assign n8584 = pi173 & ~pi221;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = ~pi173 & pi221;
  assign n8587 = ~n8585 & ~n8586;
  assign n8588 = ~n8582 & ~n8587;
  assign n8589 = ~n8581 & ~n8588;
  assign n8590 = ~n8580 & ~n8589;
  assign n8591 = ~n8579 & ~n8590;
  assign n8592 = ~n8578 & ~n8591;
  assign n8593 = ~n8577 & ~n8592;
  assign n8594 = ~n8576 & ~n8593;
  assign n8595 = ~pi169 & pi217;
  assign n8596 = ~pi168 & pi216;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = ~n8594 & n8597;
  assign n8599 = pi167 & ~pi215;
  assign n8600 = pi168 & ~pi216;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = ~n8598 & n8601;
  assign n8603 = ~n8575 & ~n8602;
  assign n8604 = ~n8574 & ~n8603;
  assign n8605 = ~pi167 & pi271;
  assign n8606 = pi169 & ~pi273;
  assign n8607 = ~pi170 & pi274;
  assign n8608 = pi170 & ~pi274;
  assign n8609 = ~pi171 & pi275;
  assign n8610 = pi171 & ~pi275;
  assign n8611 = ~pi172 & pi276;
  assign n8612 = pi172 & ~pi276;
  assign n8613 = pi174 & ~pi278;
  assign n8614 = pi173 & ~pi277;
  assign n8615 = ~n8613 & ~n8614;
  assign n8616 = ~pi173 & pi277;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = ~n8612 & ~n8617;
  assign n8619 = ~n8611 & ~n8618;
  assign n8620 = ~n8610 & ~n8619;
  assign n8621 = ~n8609 & ~n8620;
  assign n8622 = ~n8608 & ~n8621;
  assign n8623 = ~n8607 & ~n8622;
  assign n8624 = ~n8606 & ~n8623;
  assign n8625 = ~pi169 & pi273;
  assign n8626 = ~pi168 & pi272;
  assign n8627 = ~n8625 & ~n8626;
  assign n8628 = ~n8624 & n8627;
  assign n8629 = pi167 & ~pi271;
  assign n8630 = pi168 & ~pi272;
  assign n8631 = ~n8629 & ~n8630;
  assign n8632 = ~n8628 & n8631;
  assign n8633 = ~n8605 & ~n8632;
  assign n8634 = ~pi167 & pi183;
  assign n8635 = pi169 & ~pi185;
  assign n8636 = ~pi170 & pi186;
  assign n8637 = pi170 & ~pi186;
  assign n8638 = ~pi171 & pi187;
  assign n8639 = pi171 & ~pi187;
  assign n8640 = ~pi172 & pi188;
  assign n8641 = pi172 & ~pi188;
  assign n8642 = pi174 & ~pi190;
  assign n8643 = pi173 & ~pi189;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = ~pi173 & pi189;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n8641 & ~n8646;
  assign n8648 = ~n8640 & ~n8647;
  assign n8649 = ~n8639 & ~n8648;
  assign n8650 = ~n8638 & ~n8649;
  assign n8651 = ~n8637 & ~n8650;
  assign n8652 = ~n8636 & ~n8651;
  assign n8653 = ~n8635 & ~n8652;
  assign n8654 = ~pi169 & pi185;
  assign n8655 = ~pi168 & pi184;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = ~n8653 & n8656;
  assign n8658 = pi167 & ~pi183;
  assign n8659 = pi168 & ~pi184;
  assign n8660 = ~n8658 & ~n8659;
  assign n8661 = ~n8657 & n8660;
  assign n8662 = ~n8634 & ~n8661;
  assign n8663 = ~n8633 & ~n8662;
  assign n8664 = n8604 & n8663;
  assign n8665 = n8545 & n8664;
  assign n8666 = ~n8426 & n8665;
  assign n8667 = ~n3312 & ~n3678;
  assign n8668 = n6705 & n8667;
  assign n8669 = ~n2691 & ~n2841;
  assign n8670 = n5734 & n8669;
  assign n8671 = n8668 & n8670;
  assign n8672 = ~n6180 & ~n6431;
  assign n8673 = ~n7277 & ~n7533;
  assign n8674 = n8672 & n8673;
  assign n8675 = ~n4369 & ~n4647;
  assign n8676 = ~n5258 & ~n5555;
  assign n8677 = n8675 & n8676;
  assign n8678 = n8674 & n8677;
  assign n8679 = n8671 & n8678;
  assign n8680 = ~n2019 & ~n2080;
  assign n8681 = n3822 & n8680;
  assign n8682 = ~n2694 & ~n2814;
  assign n8683 = ~n4342 & ~n5231;
  assign n8684 = n8682 & n8683;
  assign n8685 = ~n3256 & ~n3651;
  assign n8686 = n4849 & n8685;
  assign n8687 = n8684 & n8686;
  assign n8688 = ~n6404 & ~n7240;
  assign n8689 = ~n7506 & n8688;
  assign n8690 = n6741 & n8689;
  assign n8691 = n8687 & n8690;
  assign n8692 = ~n998 & ~n1991;
  assign n8693 = n3858 & n8692;
  assign n8694 = n6770 & n8693;
  assign n8695 = n3942 & n5718;
  assign n8696 = n8694 & n8695;
  assign n8697 = n8691 & n8696;
  assign n8698 = ~n1172 & n8697;
  assign n8699 = ~n1025 & n8698;
  assign n8700 = ~n996 & n8699;
  assign n8701 = ~n2306 & ~n2391;
  assign n8702 = n8700 & n8701;
  assign n8703 = n3821 & n8702;
  assign n8704 = n8681 & n8703;
  assign n8705 = ~pi167 & pi175;
  assign n8706 = pi169 & ~pi177;
  assign n8707 = ~pi170 & pi178;
  assign n8708 = pi170 & ~pi178;
  assign n8709 = ~pi171 & pi179;
  assign n8710 = pi171 & ~pi179;
  assign n8711 = ~pi172 & pi180;
  assign n8712 = pi172 & ~pi180;
  assign n8713 = pi174 & ~pi182;
  assign n8714 = pi173 & ~pi181;
  assign n8715 = ~n8713 & ~n8714;
  assign n8716 = ~pi173 & pi181;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = ~n8712 & ~n8717;
  assign n8719 = ~n8711 & ~n8718;
  assign n8720 = ~n8710 & ~n8719;
  assign n8721 = ~n8709 & ~n8720;
  assign n8722 = ~n8708 & ~n8721;
  assign n8723 = ~n8707 & ~n8722;
  assign n8724 = ~n8706 & ~n8723;
  assign n8725 = ~pi169 & pi177;
  assign n8726 = ~pi168 & pi176;
  assign n8727 = ~n8725 & ~n8726;
  assign n8728 = ~n8724 & n8727;
  assign n8729 = pi167 & ~pi175;
  assign n8730 = pi168 & ~pi176;
  assign n8731 = ~n8729 & ~n8730;
  assign n8732 = ~n8728 & n8731;
  assign n8733 = ~n8705 & ~n8732;
  assign n8734 = ~pi167 & pi223;
  assign n8735 = pi169 & ~pi225;
  assign n8736 = ~pi170 & pi226;
  assign n8737 = pi170 & ~pi226;
  assign n8738 = ~pi171 & pi227;
  assign n8739 = pi171 & ~pi227;
  assign n8740 = ~pi172 & pi228;
  assign n8741 = pi172 & ~pi228;
  assign n8742 = pi174 & ~pi230;
  assign n8743 = pi173 & ~pi229;
  assign n8744 = ~n8742 & ~n8743;
  assign n8745 = ~pi173 & pi229;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = ~n8741 & ~n8746;
  assign n8748 = ~n8740 & ~n8747;
  assign n8749 = ~n8739 & ~n8748;
  assign n8750 = ~n8738 & ~n8749;
  assign n8751 = ~n8737 & ~n8750;
  assign n8752 = ~n8736 & ~n8751;
  assign n8753 = ~n8735 & ~n8752;
  assign n8754 = ~pi169 & pi225;
  assign n8755 = ~pi168 & pi224;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = ~n8753 & n8756;
  assign n8758 = pi167 & ~pi223;
  assign n8759 = pi168 & ~pi224;
  assign n8760 = ~n8758 & ~n8759;
  assign n8761 = ~n8757 & n8760;
  assign n8762 = ~n8734 & ~n8761;
  assign n8763 = ~n8733 & ~n8762;
  assign n8764 = ~pi167 & pi207;
  assign n8765 = pi169 & ~pi209;
  assign n8766 = ~pi170 & pi210;
  assign n8767 = pi170 & ~pi210;
  assign n8768 = ~pi171 & pi211;
  assign n8769 = pi171 & ~pi211;
  assign n8770 = ~pi172 & pi212;
  assign n8771 = pi172 & ~pi212;
  assign n8772 = pi174 & ~pi214;
  assign n8773 = pi173 & ~pi213;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = ~pi173 & pi213;
  assign n8776 = ~n8774 & ~n8775;
  assign n8777 = ~n8771 & ~n8776;
  assign n8778 = ~n8770 & ~n8777;
  assign n8779 = ~n8769 & ~n8778;
  assign n8780 = ~n8768 & ~n8779;
  assign n8781 = ~n8767 & ~n8780;
  assign n8782 = ~n8766 & ~n8781;
  assign n8783 = ~n8765 & ~n8782;
  assign n8784 = ~pi169 & pi209;
  assign n8785 = ~pi168 & pi208;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~n8783 & n8786;
  assign n8788 = pi167 & ~pi207;
  assign n8789 = pi168 & ~pi208;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = ~n8787 & n8790;
  assign n8792 = ~n8764 & ~n8791;
  assign n8793 = ~pi167 & pi199;
  assign n8794 = pi169 & ~pi201;
  assign n8795 = ~pi170 & pi202;
  assign n8796 = pi170 & ~pi202;
  assign n8797 = ~pi171 & pi203;
  assign n8798 = pi171 & ~pi203;
  assign n8799 = ~pi172 & pi204;
  assign n8800 = pi172 & ~pi204;
  assign n8801 = pi174 & ~pi206;
  assign n8802 = pi173 & ~pi205;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~pi173 & pi205;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = ~n8800 & ~n8805;
  assign n8807 = ~n8799 & ~n8806;
  assign n8808 = ~n8798 & ~n8807;
  assign n8809 = ~n8797 & ~n8808;
  assign n8810 = ~n8796 & ~n8809;
  assign n8811 = ~n8795 & ~n8810;
  assign n8812 = ~n8794 & ~n8811;
  assign n8813 = ~pi169 & pi201;
  assign n8814 = ~pi168 & pi200;
  assign n8815 = ~n8813 & ~n8814;
  assign n8816 = ~n8812 & n8815;
  assign n8817 = pi167 & ~pi199;
  assign n8818 = pi168 & ~pi200;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~n8816 & n8819;
  assign n8821 = ~n8793 & ~n8820;
  assign n8822 = ~n8792 & ~n8821;
  assign n8823 = n8763 & n8822;
  assign n8824 = n4787 & n8823;
  assign n8825 = n8704 & n8824;
  assign n8826 = n8679 & n8825;
  assign n8827 = n8666 & n8826;
  assign n8828 = ~n7236 & n8827;
  assign n8829 = ~n6137 & n8828;
  assign n8830 = n6193 & n8829;
  assign n8831 = n6134 & n8830;
  assign n8832 = ~n7235 & n8831;
  assign n8833 = n7296 & n8832;
  assign n8834 = n7231 & n8833;
  assign n8835 = ~n3165 & ~n3940;
  assign n8836 = ~n4001 & n8835;
  assign n8837 = ~n5043 & n8836;
  assign n8838 = ~n5943 & n8837;
  assign n8839 = ~n6951 & n8838;
  assign n8840 = ~n2934 & ~n3066;
  assign n8841 = ~n3983 & n8840;
  assign n8842 = ~n4024 & n8841;
  assign n8843 = ~n4999 & n8842;
  assign n8844 = ~n5827 & n8843;
  assign n8845 = ~n6893 & n8844;
  assign n8846 = ~n8839 & ~n8845;
  assign n8847 = ~n1086 & ~n1372;
  assign n8848 = ~n2243 & n8847;
  assign n8849 = ~n3104 & n8848;
  assign n8850 = ~n3971 & n8849;
  assign n8851 = ~n4872 & n8850;
  assign n8852 = ~n5801 & n8851;
  assign n8853 = ~n6739 & n8852;
  assign n8854 = ~n7807 & n8853;
  assign n8855 = ~n1958 & ~n2242;
  assign n8856 = ~n3095 & n8855;
  assign n8857 = ~n3997 & n8856;
  assign n8858 = ~n4837 & n8857;
  assign n8859 = ~n5822 & n8858;
  assign n8860 = ~n6820 & n8859;
  assign n8861 = ~n7785 & n8860;
  assign n8862 = ~n8854 & ~n8861;
  assign n8863 = n8846 & n8862;
  assign n8864 = ~n5469 & ~n5808;
  assign n8865 = ~n6056 & n8864;
  assign n8866 = ~n7073 & n8865;
  assign n8867 = ~n7566 & ~n7869;
  assign n8868 = ~n7240 & ~n8705;
  assign n8869 = n6740 & n8868;
  assign n8870 = n7816 & n8869;
  assign n8871 = n7814 & n8870;
  assign n8872 = n7811 & n8871;
  assign n8873 = ~n1172 & n8872;
  assign n8874 = ~n996 & n8873;
  assign n8875 = ~n2306 & n8874;
  assign n8876 = ~n500 & n8875;
  assign n8877 = n6677 & n8876;
  assign n8878 = ~n7277 & ~n8732;
  assign n8879 = n6181 & n8878;
  assign n8880 = n7279 & n8879;
  assign n8881 = n8877 & n8880;
  assign n8882 = n7284 & n8881;
  assign n8883 = ~n7236 & n8882;
  assign n8884 = ~n6137 & n8883;
  assign n8885 = n6193 & n8884;
  assign n8886 = n6134 & n8885;
  assign n8887 = ~n8867 & n8886;
  assign n8888 = ~n7235 & n8887;
  assign n8889 = n7296 & n8888;
  assign n8890 = n7231 & n8889;
  assign n8891 = ~n8866 & n8890;
  assign n8892 = ~n4163 & ~n4817;
  assign n8893 = ~n4902 & n8892;
  assign n8894 = ~n6001 & n8893;
  assign n8895 = ~n7014 & n8894;
  assign n8896 = ~n6282 & ~n6784;
  assign n8897 = ~n7158 & n8896;
  assign n8898 = ~n8895 & ~n8897;
  assign n8899 = n8891 & n8898;
  assign n8900 = n8863 & n8899;
  assign n8901 = ~n8834 & ~n8900;
  assign po165 = n8397 | ~n8901;
  assign n8903 = ~n8378 & ~po165;
  assign n8904 = pi016 & ~n8391;
  assign n8905 = ~po161 & n8904;
  assign n8906 = ~n8017 & n8905;
  assign n8907 = ~n8314 & n8906;
  assign n8908 = n8281 & n8907;
  assign n8909 = n8390 & n8908;
  assign n8910 = n8383 & n8909;
  assign n8911 = n7241 & ~n8705;
  assign n8912 = n5724 & n8911;
  assign n8913 = pi018 & ~n501;
  assign n8914 = n5714 & n8913;
  assign n8915 = n5719 & n8914;
  assign n8916 = n8912 & n8915;
  assign n8917 = ~n1172 & n8916;
  assign n8918 = ~n996 & n8917;
  assign n8919 = ~n2306 & n8918;
  assign n8920 = ~n500 & n8919;
  assign n8921 = n6677 & n8920;
  assign n8922 = n8880 & n8921;
  assign n8923 = n7284 & n8922;
  assign n8924 = ~n7236 & n8923;
  assign n8925 = ~n6137 & n8924;
  assign n8926 = n6193 & n8925;
  assign n8927 = n6134 & n8926;
  assign n8928 = ~n8867 & n8927;
  assign n8929 = ~n7235 & n8928;
  assign n8930 = n7296 & n8929;
  assign n8931 = n7231 & n8930;
  assign n8932 = ~n8866 & n8931;
  assign n8933 = n8898 & n8932;
  assign n8934 = n8863 & n8933;
  assign n8935 = n5720 & n8685;
  assign n8936 = n4797 & n8935;
  assign n8937 = ~n6404 & ~n7506;
  assign n8938 = n7241 & n8937;
  assign n8939 = n8684 & n8938;
  assign n8940 = n8936 & n8939;
  assign n8941 = n4792 & n5754;
  assign n8942 = pi017 & ~n501;
  assign n8943 = n8692 & n8942;
  assign n8944 = n8941 & n8943;
  assign n8945 = n3810 & n5717;
  assign n8946 = n4790 & n8945;
  assign n8947 = n8944 & n8946;
  assign n8948 = n8940 & n8947;
  assign n8949 = ~n1172 & n8948;
  assign n8950 = ~n1025 & n8949;
  assign n8951 = ~n996 & n8950;
  assign n8952 = n8701 & n8951;
  assign n8953 = n3821 & n8952;
  assign n8954 = n8681 & n8953;
  assign n8955 = n8824 & n8954;
  assign n8956 = n8679 & n8955;
  assign n8957 = n8666 & n8956;
  assign n8958 = ~n7236 & n8957;
  assign n8959 = ~n6137 & n8958;
  assign n8960 = n6193 & n8959;
  assign n8961 = n6134 & n8960;
  assign n8962 = ~n7235 & n8961;
  assign n8963 = n7296 & n8962;
  assign n8964 = n7231 & n8963;
  assign n8965 = ~n8934 & ~n8964;
  assign n8966 = ~n8910 & n8965;
  assign po009 = n8903 | ~n8966;
  assign n8968 = n7898 & ~n8397;
  assign n8969 = ~n1026 & ~n1115;
  assign n8970 = ~n1086 & n8969;
  assign n8971 = ~n1208 & n8970;
  assign n8972 = n4920 & n8971;
  assign n8973 = ~n1270 & n8972;
  assign n8974 = n4932 & n8973;
  assign n8975 = ~n1372 & n8974;
  assign n8976 = ~n2243 & n8975;
  assign n8977 = ~n3104 & n8976;
  assign n8978 = ~n3837 & n8977;
  assign n8979 = ~n3971 & n8978;
  assign n8980 = ~n4872 & n8979;
  assign n8981 = ~n5801 & n8980;
  assign n8982 = ~n6739 & n8981;
  assign n8983 = ~n7945 & n8982;
  assign n8984 = ~n7944 & n8983;
  assign n8985 = ~n7807 & n8984;
  assign n8986 = ~n7943 & n8985;
  assign n8987 = n7966 & n8986;
  assign n8988 = n7942 & n8987;
  assign n8989 = n7935 & n8988;
  assign n8990 = n7895 & ~n8989;
  assign n8991 = ~n8968 & ~n8990;
  assign n8992 = n7924 & ~n8250;
  assign n8993 = n7894 & ~n8291;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = n8991 & n8994;
  assign n8996 = n7905 & ~n8037;
  assign n8997 = ~n7890 & n7892;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = n7923 & ~n8114;
  assign n9000 = n7907 & ~n8346;
  assign n9001 = ~n8999 & ~n9000;
  assign n9002 = n8998 & n9001;
  assign n9003 = n7901 & ~n8053;
  assign n9004 = n7902 & ~n8218;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = n1958 & ~n8900;
  assign n9007 = n7899 & ~n8145;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = n9005 & n9008;
  assign n9010 = n7891 & ~n8179;
  assign n9011 = ~n1897 & ~n1958;
  assign n9012 = n4828 & n9011;
  assign n9013 = n1743 & n9012;
  assign n9014 = ~n2242 & n9013;
  assign n9015 = ~n3095 & n9014;
  assign n9016 = ~n3997 & n9015;
  assign n9017 = ~n4003 & n9016;
  assign n9018 = ~n4837 & n9017;
  assign n9019 = ~n5822 & n9018;
  assign n9020 = ~n6820 & n9019;
  assign n9021 = ~n7907 & n9020;
  assign n9022 = ~n7906 & n9021;
  assign n9023 = ~n7785 & n9022;
  assign n9024 = ~n7905 & n9023;
  assign n9025 = n7925 & n9024;
  assign n9026 = n7904 & n9025;
  assign n9027 = n7897 & n9026;
  assign n9028 = n7906 & ~n7999;
  assign n9029 = n2020 & ~n8834;
  assign n9030 = ~n1897 & n2255;
  assign n9031 = n1743 & n9030;
  assign n9032 = ~n2242 & n9031;
  assign n9033 = ~n3095 & n9032;
  assign n9034 = ~n3997 & n9033;
  assign n9035 = ~n4003 & n9034;
  assign n9036 = ~n4837 & n9035;
  assign n9037 = ~n5822 & n9036;
  assign n9038 = ~n6820 & n9037;
  assign n9039 = ~n7785 & n9038;
  assign n9040 = ~n9029 & n9039;
  assign n9041 = ~n9028 & n9040;
  assign n9042 = ~n9027 & n9041;
  assign n9043 = ~n9010 & n9042;
  assign n9044 = n9009 & n9043;
  assign n9045 = n9002 & n9044;
  assign n9046 = n8995 & n9045;
  assign n9047 = n7965 & ~n8037;
  assign n9048 = ~n7890 & n7943;
  assign n9049 = ~n9047 & ~n9048;
  assign n9050 = n7929 & ~n8114;
  assign n9051 = n7964 & ~n8291;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = n9049 & n9052;
  assign n9054 = n7936 & ~n8397;
  assign n9055 = n7933 & ~n9027;
  assign n9056 = ~n9054 & ~n9055;
  assign n9057 = n7930 & ~n8250;
  assign n9058 = n7932 & ~n8179;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = n9056 & n9059;
  assign n9061 = n7940 & ~n8218;
  assign n9062 = n1086 & ~n8900;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = n7937 & ~n8145;
  assign n9065 = ~n8989 & ~n9064;
  assign n9066 = n9063 & n9065;
  assign n9067 = n7945 & ~n8346;
  assign n9068 = n7939 & ~n8053;
  assign n9069 = n7944 & ~n7999;
  assign n9070 = n1026 & ~n8834;
  assign n9071 = ~n1208 & n7946;
  assign n9072 = n4920 & n9071;
  assign n9073 = ~n1270 & n9072;
  assign n9074 = n4932 & n9073;
  assign n9075 = ~n1372 & n9074;
  assign n9076 = ~n2243 & n9075;
  assign n9077 = ~n3104 & n9076;
  assign n9078 = ~n3971 & n9077;
  assign n9079 = ~n4003 & n9078;
  assign n9080 = ~n4872 & n9079;
  assign n9081 = ~n5801 & n9080;
  assign n9082 = ~n6739 & n9081;
  assign n9083 = ~n7807 & n9082;
  assign n9084 = ~n9070 & n9083;
  assign n9085 = ~n9069 & n9084;
  assign n9086 = ~n9068 & n9085;
  assign n9087 = ~n9067 & n9086;
  assign n9088 = n9066 & n9087;
  assign n9089 = n9060 & n9088;
  assign n9090 = n9053 & n9089;
  assign n9091 = n7834 & ~n8397;
  assign n9092 = n7808 & ~n8989;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = n7786 & ~n9027;
  assign n9095 = n7788 & ~n8291;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = n9093 & n9096;
  assign n9098 = n7885 & ~n8114;
  assign n9099 = n7841 & ~n8037;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = n7767 & ~n8179;
  assign n9102 = n7886 & ~n8250;
  assign n9103 = ~n9101 & ~n9102;
  assign n9104 = n9100 & n9103;
  assign n9105 = n7837 & ~n8053;
  assign n9106 = n7838 & ~n8218;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = n2934 & ~n8900;
  assign n9109 = n7835 & ~n8145;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = n9107 & n9110;
  assign n9112 = n7870 & ~n8346;
  assign n9113 = n7842 & ~n7999;
  assign n9114 = n2842 & ~n8834;
  assign n9115 = ~n2663 & n2784;
  assign n9116 = ~n3024 & n9115;
  assign n9117 = n2634 & n9116;
  assign n9118 = ~n3066 & n9117;
  assign n9119 = ~n3983 & n9118;
  assign n9120 = ~n4003 & n9119;
  assign n9121 = ~n4024 & n9120;
  assign n9122 = ~n4999 & n9121;
  assign n9123 = ~n5827 & n9122;
  assign n9124 = ~n6893 & n9123;
  assign n9125 = ~n9114 & n9124;
  assign n9126 = ~n9113 & n9125;
  assign n9127 = ~n7890 & n9126;
  assign n9128 = ~n9112 & n9127;
  assign n9129 = n9111 & n9128;
  assign n9130 = n9104 & n9129;
  assign n9131 = n9097 & n9130;
  assign n9132 = ~n9090 & ~n9131;
  assign n9133 = ~n9046 & n9132;
  assign n9134 = n3846 & n7972;
  assign n9135 = n3854 & n9134;
  assign n9136 = ~n2663 & ~n2783;
  assign n9137 = n3849 & n9136;
  assign n9138 = ~n3024 & n9137;
  assign n9139 = n9135 & n9138;
  assign n9140 = ~n3066 & n9139;
  assign n9141 = ~n3983 & n9140;
  assign n9142 = ~n4003 & n9141;
  assign n9143 = ~n4024 & n9142;
  assign n9144 = ~n4999 & n9143;
  assign n9145 = ~n5827 & n9144;
  assign n9146 = ~n6893 & n9145;
  assign n9147 = ~n9114 & n9146;
  assign n9148 = ~n9113 & n9147;
  assign n9149 = ~n7890 & n9148;
  assign n9150 = ~n9112 & n9149;
  assign n9151 = n9111 & n9150;
  assign n9152 = n9104 & n9151;
  assign n9153 = n9097 & n9152;
  assign n9154 = ~n7890 & n7997;
  assign n9155 = n7994 & ~n7999;
  assign n9156 = ~n9154 & n9155;
  assign n9157 = n7993 & ~n9027;
  assign n9158 = n7996 & ~n8989;
  assign n9159 = ~n9157 & ~n9158;
  assign n9160 = n9156 & n9159;
  assign n9161 = ~n9153 & ~n9160;
  assign n9162 = ~n9133 & n9161;
  assign n9163 = n8009 & ~n8397;
  assign n9164 = n8006 & ~n8989;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = n8018 & ~n8346;
  assign n9167 = n8032 & ~n8291;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = n9165 & n9168;
  assign n9170 = n8016 & ~n8114;
  assign n9171 = ~n7890 & n8003;
  assign n9172 = ~n9170 & ~n9171;
  assign n9173 = n8033 & ~n8179;
  assign n9174 = n8005 & ~n9027;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = n9172 & n9175;
  assign n9177 = n8012 & ~n8053;
  assign n9178 = n8013 & ~n8218;
  assign n9179 = ~n9177 & ~n9178;
  assign n9180 = n3165 & ~n8900;
  assign n9181 = n8010 & ~n8145;
  assign n9182 = ~n9180 & ~n9181;
  assign n9183 = n9179 & n9182;
  assign n9184 = n8002 & ~n8250;
  assign n9185 = ~n7999 & n8017;
  assign n9186 = n3679 & ~n8834;
  assign n9187 = ~n3464 & n8056;
  assign n9188 = n8020 & n9187;
  assign n9189 = ~n3940 & n9188;
  assign n9190 = ~n4001 & n9189;
  assign n9191 = ~n5043 & n9190;
  assign n9192 = ~n5943 & n9191;
  assign n9193 = ~n6951 & n9192;
  assign n9194 = ~n9186 & n9193;
  assign n9195 = ~n9185 & n9194;
  assign n9196 = ~n8037 & n9195;
  assign n9197 = ~n9184 & n9196;
  assign n9198 = n9183 & n9197;
  assign n9199 = n9176 & n9198;
  assign n9200 = n9169 & n9199;
  assign n9201 = ~n7999 & n8039;
  assign n9202 = ~n9154 & n9201;
  assign n9203 = n9159 & n9202;
  assign n9204 = ~n9200 & ~n9203;
  assign n9205 = ~n9162 & n9204;
  assign n9206 = n8050 & ~n8989;
  assign n9207 = n8045 & ~n8053;
  assign n9208 = ~n9185 & n9207;
  assign n9209 = ~n9206 & n9208;
  assign n9210 = ~n8037 & n8049;
  assign n9211 = ~n7890 & n8044;
  assign n9212 = n8048 & ~n9027;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9210 & n9213;
  assign n9215 = n9209 & n9214;
  assign n9216 = n3740 & n8054;
  assign n9217 = n3951 & n9216;
  assign n9218 = ~n3344 & ~n3650;
  assign n9219 = n4100 & n9218;
  assign n9220 = ~n3464 & n9219;
  assign n9221 = n9217 & n9220;
  assign n9222 = ~n3940 & n9221;
  assign n9223 = ~n4001 & n9222;
  assign n9224 = ~n5043 & n9223;
  assign n9225 = ~n5943 & n9224;
  assign n9226 = ~n6951 & n9225;
  assign n9227 = ~n9186 & n9226;
  assign n9228 = ~n9185 & n9227;
  assign n9229 = ~n8037 & n9228;
  assign n9230 = ~n9184 & n9229;
  assign n9231 = n9183 & n9230;
  assign n9232 = n9176 & n9231;
  assign n9233 = n9169 & n9232;
  assign n9234 = ~n9215 & ~n9233;
  assign n9235 = ~n9205 & n9234;
  assign n9236 = ~n8053 & n8076;
  assign n9237 = ~n9185 & n9236;
  assign n9238 = ~n9206 & n9237;
  assign n9239 = n9214 & n9238;
  assign n9240 = ~n8037 & n8080;
  assign n9241 = ~n7890 & n8081;
  assign n9242 = ~n9240 & ~n9241;
  assign n9243 = n8093 & ~n8179;
  assign n9244 = n8109 & ~n8291;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = n9242 & n9245;
  assign n9247 = n8090 & ~n8397;
  assign n9248 = n8084 & ~n8989;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = n8094 & ~n8346;
  assign n9251 = n8110 & ~n8250;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = n9249 & n9252;
  assign n9254 = n8087 & ~n8218;
  assign n9255 = ~n9207 & ~n9254;
  assign n9256 = n4163 & ~n8900;
  assign n9257 = n8089 & ~n8145;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = n9255 & n9258;
  assign n9260 = n8083 & ~n9027;
  assign n9261 = n4370 & ~n8834;
  assign n9262 = ~n4341 & ~n4579;
  assign n9263 = ~n4608 & n9262;
  assign n9264 = ~n4192 & n9263;
  assign n9265 = n8098 & n9264;
  assign n9266 = ~n4817 & n9265;
  assign n9267 = ~n4902 & n9266;
  assign n9268 = ~n6001 & n9267;
  assign n9269 = ~n7014 & n9268;
  assign n9270 = ~n9261 & n9269;
  assign n9271 = ~n9185 & n9270;
  assign n9272 = ~n8114 & n9271;
  assign n9273 = ~n9260 & n9272;
  assign n9274 = n9259 & n9273;
  assign n9275 = n9253 & n9274;
  assign n9276 = n9246 & n9275;
  assign n9277 = ~n9239 & ~n9276;
  assign n9278 = ~n9235 & n9277;
  assign n9279 = n4737 & n8117;
  assign n9280 = n4491 & n9279;
  assign n9281 = n4609 & n5094;
  assign n9282 = ~n4192 & n9281;
  assign n9283 = n9280 & n9282;
  assign n9284 = ~n4817 & n9283;
  assign n9285 = ~n4902 & n9284;
  assign n9286 = ~n6001 & n9285;
  assign n9287 = ~n7014 & n9286;
  assign n9288 = ~n9261 & n9287;
  assign n9289 = ~n9185 & n9288;
  assign n9290 = ~n8114 & n9289;
  assign n9291 = ~n9260 & n9290;
  assign n9292 = n9259 & n9291;
  assign n9293 = n9253 & n9292;
  assign n9294 = n9246 & n9293;
  assign n9295 = n8135 & ~n8989;
  assign n9296 = ~n7890 & n8133;
  assign n9297 = n8142 & ~n9027;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = ~n9295 & n9298;
  assign n9300 = n8138 & ~n8145;
  assign n9301 = ~n9185 & n9300;
  assign n9302 = ~n9207 & n9301;
  assign n9303 = ~n8037 & n8134;
  assign n9304 = ~n8114 & n8141;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = n9302 & n9305;
  assign n9307 = n9299 & n9306;
  assign n9308 = ~n9294 & ~n9307;
  assign n9309 = ~n9278 & n9308;
  assign n9310 = ~n8037 & n8175;
  assign n9311 = ~n7890 & n8149;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = ~n8114 & n8160;
  assign n9314 = n8174 & ~n8291;
  assign n9315 = ~n9313 & ~n9314;
  assign n9316 = n9312 & n9315;
  assign n9317 = n8156 & ~n8397;
  assign n9318 = n8151 & ~n8989;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = n8161 & ~n8346;
  assign n9321 = n8148 & ~n8250;
  assign n9322 = ~n9320 & ~n9321;
  assign n9323 = n9319 & n9322;
  assign n9324 = ~n9207 & ~n9300;
  assign n9325 = n8157 & ~n8218;
  assign n9326 = n5469 & ~n8900;
  assign n9327 = ~n9325 & ~n9326;
  assign n9328 = n9324 & n9327;
  assign n9329 = n8152 & ~n9027;
  assign n9330 = n5259 & ~n8834;
  assign n9331 = ~n5230 & ~n5289;
  assign n9332 = ~n5527 & n9331;
  assign n9333 = ~n5170 & n9332;
  assign n9334 = n8162 & n9333;
  assign n9335 = ~n5808 & n9334;
  assign n9336 = ~n6056 & n9335;
  assign n9337 = ~n7073 & n9336;
  assign n9338 = ~n9330 & n9337;
  assign n9339 = ~n9185 & n9338;
  assign n9340 = ~n8179 & n9339;
  assign n9341 = ~n9329 & n9340;
  assign n9342 = n9328 & n9341;
  assign n9343 = n9323 & n9342;
  assign n9344 = n9316 & n9343;
  assign n9345 = ~n8145 & n8182;
  assign n9346 = ~n9185 & n9345;
  assign n9347 = ~n9207 & n9346;
  assign n9348 = n9305 & n9347;
  assign n9349 = n9299 & n9348;
  assign n9350 = ~n9344 & ~n9349;
  assign n9351 = ~n9309 & n9350;
  assign n9352 = n6068 & n8189;
  assign n9353 = n6066 & n9352;
  assign n9354 = n6073 & n8163;
  assign n9355 = ~n5170 & n9354;
  assign n9356 = n9353 & n9355;
  assign n9357 = ~n5808 & n9356;
  assign n9358 = ~n6056 & n9357;
  assign n9359 = ~n7073 & n9358;
  assign n9360 = ~n9330 & n9359;
  assign n9361 = ~n9185 & n9360;
  assign n9362 = ~n8179 & n9361;
  assign n9363 = ~n9329 & n9362;
  assign n9364 = n9328 & n9363;
  assign n9365 = n9323 & n9364;
  assign n9366 = n9316 & n9365;
  assign n9367 = ~n7890 & n8207;
  assign n9368 = ~n8114 & n8215;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = n8208 & ~n8989;
  assign n9371 = n8214 & ~n9027;
  assign n9372 = ~n9370 & ~n9371;
  assign n9373 = n9369 & n9372;
  assign n9374 = n8211 & ~n8218;
  assign n9375 = ~n9185 & n9374;
  assign n9376 = n9324 & n9375;
  assign n9377 = ~n8179 & n8205;
  assign n9378 = ~n8037 & n8204;
  assign n9379 = ~n9377 & ~n9378;
  assign n9380 = n9376 & n9379;
  assign n9381 = n9373 & n9380;
  assign n9382 = ~n9366 & ~n9381;
  assign n9383 = ~n9351 & n9382;
  assign n9384 = ~n8037 & n8231;
  assign n9385 = ~n7890 & n8221;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = ~n8114 & n8245;
  assign n9388 = n8224 & ~n8291;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = n9386 & n9389;
  assign n9391 = n8228 & ~n8397;
  assign n9392 = n8246 & ~n8989;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = n8232 & ~n8346;
  assign n9395 = ~n8179 & n8222;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = n9393 & n9396;
  assign n9398 = n6282 & ~n8900;
  assign n9399 = ~n9374 & ~n9398;
  assign n9400 = n9324 & n9399;
  assign n9401 = n8225 & ~n9027;
  assign n9402 = n6432 & ~n8834;
  assign n9403 = n7170 & n7177;
  assign n9404 = ~n6224 & n8261;
  assign n9405 = n9403 & n9404;
  assign n9406 = ~n6784 & n9405;
  assign n9407 = ~n7158 & n9406;
  assign n9408 = ~n9402 & n9407;
  assign n9409 = ~n9185 & n9408;
  assign n9410 = ~n8250 & n9409;
  assign n9411 = ~n9401 & n9410;
  assign n9412 = n9400 & n9411;
  assign n9413 = n9397 & n9412;
  assign n9414 = n9390 & n9413;
  assign n9415 = ~n8218 & n8252;
  assign n9416 = ~n9185 & n9415;
  assign n9417 = n9324 & n9416;
  assign n9418 = n9379 & n9417;
  assign n9419 = n9373 & n9418;
  assign n9420 = ~n9414 & ~n9419;
  assign n9421 = ~n9383 & n9420;
  assign n9422 = ~pi013 & ~n6461;
  assign n9423 = n6343 & n9422;
  assign n9424 = n8233 & n9423;
  assign n9425 = ~n6224 & n8236;
  assign n9426 = n9424 & n9425;
  assign n9427 = ~n6784 & n9426;
  assign n9428 = ~n7158 & n9427;
  assign n9429 = ~n9402 & n9428;
  assign n9430 = ~n9185 & n9429;
  assign n9431 = ~n8250 & n9430;
  assign n9432 = ~n9401 & n9431;
  assign n9433 = n9400 & n9432;
  assign n9434 = n9397 & n9433;
  assign n9435 = n9390 & n9434;
  assign n9436 = ~n8250 & n8277;
  assign n9437 = ~n8179 & n8278;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = ~n7890 & n8274;
  assign n9440 = ~n8114 & n8275;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = n9438 & n9441;
  assign n9443 = n9324 & ~n9374;
  assign n9444 = n8286 & ~n8989;
  assign n9445 = n8314 & ~n9185;
  assign n9446 = ~n8291 & n9445;
  assign n9447 = ~n9444 & n9446;
  assign n9448 = n8287 & ~n9027;
  assign n9449 = ~n8037 & n8282;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = n9447 & n9450;
  assign n9452 = n9443 & n9451;
  assign n9453 = n9442 & n9452;
  assign n9454 = ~n8037 & n8304;
  assign n9455 = ~n7890 & n8297;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = ~n8114 & n8335;
  assign n9458 = ~n8291 & n8314;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = n9456 & n9459;
  assign n9461 = n8329 & ~n8397;
  assign n9462 = n8323 & ~n8989;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = ~n8250 & n8299;
  assign n9465 = ~n8179 & n8326;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = n9463 & n9466;
  assign n9468 = n7566 & ~n8900;
  assign n9469 = ~n9374 & ~n9468;
  assign n9470 = n9324 & n9469;
  assign n9471 = n8313 & ~n9027;
  assign n9472 = n7534 & ~n8834;
  assign n9473 = ~n7327 & ~n7505;
  assign n9474 = n7476 & n9473;
  assign n9475 = n7753 & n9474;
  assign n9476 = ~n7595 & n8363;
  assign n9477 = n9475 & n9476;
  assign n9478 = ~n7869 & n9477;
  assign n9479 = ~n9472 & n9478;
  assign n9480 = ~n9185 & n9479;
  assign n9481 = ~n8346 & n9480;
  assign n9482 = ~n9471 & n9481;
  assign n9483 = n9470 & n9482;
  assign n9484 = n9467 & n9483;
  assign n9485 = n9460 & n9484;
  assign n9486 = ~n9453 & ~n9485;
  assign n9487 = ~n9435 & n9486;
  assign n9488 = ~n9421 & n9487;
  assign n9489 = ~n7204 & n8350;
  assign n9490 = ~n9185 & n9489;
  assign n9491 = ~n8291 & n9490;
  assign n9492 = ~n9444 & n9491;
  assign n9493 = n9450 & n9492;
  assign n9494 = n9443 & n9493;
  assign n9495 = n9442 & n9494;
  assign n9496 = n8359 & n8364;
  assign n9497 = n8357 & n8358;
  assign n9498 = n9496 & n9497;
  assign n9499 = n7417 & ~n7595;
  assign n9500 = n9498 & n9499;
  assign n9501 = ~n7869 & n9500;
  assign n9502 = ~n9472 & n9501;
  assign n9503 = ~n9185 & n9502;
  assign n9504 = ~n8346 & n9503;
  assign n9505 = ~n9471 & n9504;
  assign n9506 = n9470 & n9505;
  assign n9507 = n9467 & n9506;
  assign n9508 = n9460 & n9507;
  assign n9509 = ~n9495 & ~n9508;
  assign n9510 = ~n9488 & n9509;
  assign n9511 = ~n8733 & ~n8834;
  assign n9512 = ~n8900 & ~n9511;
  assign n9513 = ~n9185 & n9512;
  assign n9514 = ~n9458 & n9513;
  assign n9515 = ~po161 & ~n8397;
  assign n9516 = n8861 & ~n9027;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = n9514 & n9517;
  assign n9519 = n9443 & n9518;
  assign n9520 = ~n8114 & n8895;
  assign n9521 = ~n8179 & n8866;
  assign n9522 = ~n8037 & n8839;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = ~n9520 & n9523;
  assign n9525 = ~n8346 & n8867;
  assign n9526 = n8854 & ~n8989;
  assign n9527 = ~n9525 & ~n9526;
  assign n9528 = ~n8250 & n8897;
  assign n9529 = ~n7890 & n8845;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = n9527 & n9530;
  assign n9532 = n9524 & n9531;
  assign n9533 = n9519 & n9532;
  assign n9534 = ~pi183 & pi207;
  assign n9535 = pi183 & ~pi207;
  assign n9536 = ~pi184 & pi208;
  assign n9537 = pi184 & ~pi208;
  assign n9538 = ~pi185 & pi209;
  assign n9539 = pi185 & ~pi209;
  assign n9540 = ~pi186 & pi210;
  assign n9541 = pi186 & ~pi210;
  assign n9542 = ~pi187 & pi211;
  assign n9543 = pi187 & ~pi211;
  assign n9544 = ~pi189 & pi213;
  assign n9545 = pi190 & ~pi214;
  assign n9546 = ~n9544 & n9545;
  assign n9547 = pi189 & ~pi213;
  assign n9548 = pi188 & ~pi212;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~n9546 & n9549;
  assign n9551 = ~pi188 & pi212;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = ~n9543 & ~n9552;
  assign n9554 = ~n9542 & ~n9553;
  assign n9555 = ~n9541 & ~n9554;
  assign n9556 = ~n9540 & ~n9555;
  assign n9557 = ~n9539 & ~n9556;
  assign n9558 = ~n9538 & ~n9557;
  assign n9559 = ~n9537 & ~n9558;
  assign n9560 = ~n9536 & ~n9559;
  assign n9561 = ~n9535 & ~n9560;
  assign n9562 = ~n9534 & ~n9561;
  assign n9563 = pi184 & ~pi200;
  assign n9564 = ~pi185 & pi201;
  assign n9565 = pi185 & ~pi201;
  assign n9566 = ~pi186 & pi202;
  assign n9567 = pi186 & ~pi202;
  assign n9568 = ~pi187 & pi203;
  assign n9569 = pi187 & ~pi203;
  assign n9570 = ~pi189 & pi205;
  assign n9571 = pi190 & ~pi206;
  assign n9572 = ~n9570 & n9571;
  assign n9573 = pi189 & ~pi205;
  assign n9574 = pi188 & ~pi204;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = ~n9572 & n9575;
  assign n9577 = ~pi188 & pi204;
  assign n9578 = ~n9576 & ~n9577;
  assign n9579 = ~n9569 & ~n9578;
  assign n9580 = ~n9568 & ~n9579;
  assign n9581 = ~n9567 & ~n9580;
  assign n9582 = ~n9566 & ~n9581;
  assign n9583 = ~n9565 & ~n9582;
  assign n9584 = ~n9564 & ~n9583;
  assign n9585 = ~n9563 & ~n9584;
  assign n9586 = ~pi184 & pi200;
  assign n9587 = pi183 & ~n9586;
  assign n9588 = ~n9585 & n9587;
  assign n9589 = pi199 & ~n9588;
  assign n9590 = ~n9585 & ~n9586;
  assign n9591 = ~pi183 & ~n9590;
  assign n9592 = ~n9589 & ~n9591;
  assign n9593 = pi184 & ~pi224;
  assign n9594 = ~pi185 & pi225;
  assign n9595 = pi185 & ~pi225;
  assign n9596 = ~pi186 & pi226;
  assign n9597 = pi186 & ~pi226;
  assign n9598 = ~pi187 & pi227;
  assign n9599 = pi187 & ~pi227;
  assign n9600 = ~pi189 & pi229;
  assign n9601 = pi190 & ~pi230;
  assign n9602 = ~n9600 & n9601;
  assign n9603 = pi189 & ~pi229;
  assign n9604 = pi188 & ~pi228;
  assign n9605 = ~n9603 & ~n9604;
  assign n9606 = ~n9602 & n9605;
  assign n9607 = ~pi188 & pi228;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~n9599 & ~n9608;
  assign n9610 = ~n9598 & ~n9609;
  assign n9611 = ~n9597 & ~n9610;
  assign n9612 = ~n9596 & ~n9611;
  assign n9613 = ~n9595 & ~n9612;
  assign n9614 = ~n9594 & ~n9613;
  assign n9615 = ~n9593 & ~n9614;
  assign n9616 = ~pi184 & pi224;
  assign n9617 = pi183 & ~n9616;
  assign n9618 = ~n9615 & n9617;
  assign n9619 = pi223 & ~n9618;
  assign n9620 = ~n9615 & ~n9616;
  assign n9621 = ~pi183 & ~n9620;
  assign n9622 = ~n9619 & ~n9621;
  assign n9623 = ~n9592 & ~n9622;
  assign n9624 = ~n9562 & n9623;
  assign n9625 = pi184 & ~pi192;
  assign n9626 = ~pi185 & pi193;
  assign n9627 = pi185 & ~pi193;
  assign n9628 = ~pi186 & pi194;
  assign n9629 = pi186 & ~pi194;
  assign n9630 = ~pi187 & pi195;
  assign n9631 = pi187 & ~pi195;
  assign n9632 = ~pi189 & pi197;
  assign n9633 = pi190 & ~pi198;
  assign n9634 = ~n9632 & n9633;
  assign n9635 = pi189 & ~pi197;
  assign n9636 = pi188 & ~pi196;
  assign n9637 = ~n9635 & ~n9636;
  assign n9638 = ~n9634 & n9637;
  assign n9639 = ~pi188 & pi196;
  assign n9640 = ~n9638 & ~n9639;
  assign n9641 = ~n9631 & ~n9640;
  assign n9642 = ~n9630 & ~n9641;
  assign n9643 = ~n9629 & ~n9642;
  assign n9644 = ~n9628 & ~n9643;
  assign n9645 = ~n9627 & ~n9644;
  assign n9646 = ~n9626 & ~n9645;
  assign n9647 = ~n9625 & ~n9646;
  assign n9648 = ~pi184 & pi192;
  assign n9649 = pi183 & ~n9648;
  assign n9650 = ~n9647 & n9649;
  assign n9651 = pi191 & ~n9650;
  assign n9652 = ~n9647 & ~n9648;
  assign n9653 = ~pi183 & ~n9652;
  assign n9654 = ~n9651 & ~n9653;
  assign n9655 = ~n7326 & ~n8661;
  assign n9656 = n8878 & n9655;
  assign n9657 = ~n9654 & n9656;
  assign n9658 = pi184 & ~pi216;
  assign n9659 = ~pi185 & pi217;
  assign n9660 = pi185 & ~pi217;
  assign n9661 = ~pi186 & pi218;
  assign n9662 = pi186 & ~pi218;
  assign n9663 = ~pi187 & pi219;
  assign n9664 = pi187 & ~pi219;
  assign n9665 = ~pi189 & pi221;
  assign n9666 = pi190 & ~pi222;
  assign n9667 = ~n9665 & n9666;
  assign n9668 = pi189 & ~pi221;
  assign n9669 = pi188 & ~pi220;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = ~n9667 & n9670;
  assign n9672 = ~pi188 & pi220;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = ~n9664 & ~n9673;
  assign n9675 = ~n9663 & ~n9674;
  assign n9676 = ~n9662 & ~n9675;
  assign n9677 = ~n9661 & ~n9676;
  assign n9678 = ~n9660 & ~n9677;
  assign n9679 = ~n9659 & ~n9678;
  assign n9680 = ~n9658 & ~n9679;
  assign n9681 = ~pi184 & pi216;
  assign n9682 = pi183 & ~n9681;
  assign n9683 = ~n9680 & n9682;
  assign n9684 = pi215 & ~n9683;
  assign n9685 = ~n9680 & ~n9681;
  assign n9686 = ~pi183 & ~n9685;
  assign n9687 = ~n9684 & ~n9686;
  assign n9688 = pi184 & ~pi232;
  assign n9689 = ~pi185 & pi233;
  assign n9690 = pi185 & ~pi233;
  assign n9691 = ~pi186 & pi234;
  assign n9692 = pi186 & ~pi234;
  assign n9693 = ~pi187 & pi235;
  assign n9694 = pi187 & ~pi235;
  assign n9695 = ~pi189 & pi237;
  assign n9696 = pi190 & ~pi238;
  assign n9697 = ~n9695 & n9696;
  assign n9698 = pi189 & ~pi237;
  assign n9699 = pi188 & ~pi236;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = ~n9697 & n9700;
  assign n9702 = ~pi188 & pi236;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = ~n9694 & ~n9703;
  assign n9705 = ~n9693 & ~n9704;
  assign n9706 = ~n9692 & ~n9705;
  assign n9707 = ~n9691 & ~n9706;
  assign n9708 = ~n9690 & ~n9707;
  assign n9709 = ~n9689 & ~n9708;
  assign n9710 = ~n9688 & ~n9709;
  assign n9711 = ~pi184 & pi232;
  assign n9712 = pi183 & ~n9711;
  assign n9713 = ~n9710 & n9712;
  assign n9714 = pi231 & ~n9713;
  assign n9715 = ~n9710 & ~n9711;
  assign n9716 = ~pi183 & ~n9715;
  assign n9717 = ~n9714 & ~n9716;
  assign n9718 = ~n9687 & ~n9717;
  assign n9719 = n9657 & n9718;
  assign n9720 = ~n3312 & ~n3523;
  assign n9721 = n5734 & n9720;
  assign n9722 = ~n2452 & ~n2691;
  assign n9723 = n8701 & n9722;
  assign n9724 = n9721 & n9723;
  assign n9725 = ~n5526 & ~n5555;
  assign n9726 = ~n6180 & ~n6460;
  assign n9727 = n9725 & n9726;
  assign n9728 = ~n4647 & ~n4676;
  assign n9729 = n6705 & n9728;
  assign n9730 = n9727 & n9729;
  assign n9731 = n9724 & n9730;
  assign n9732 = n9719 & n9731;
  assign n9733 = n9624 & n9732;
  assign n9734 = pi184 & ~pi272;
  assign n9735 = ~pi185 & pi273;
  assign n9736 = pi185 & ~pi273;
  assign n9737 = ~pi186 & pi274;
  assign n9738 = pi186 & ~pi274;
  assign n9739 = ~pi187 & pi275;
  assign n9740 = pi187 & ~pi275;
  assign n9741 = ~pi188 & pi276;
  assign n9742 = pi188 & ~pi276;
  assign n9743 = pi190 & ~pi278;
  assign n9744 = pi189 & ~pi277;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = ~pi189 & pi277;
  assign n9747 = ~n9745 & ~n9746;
  assign n9748 = ~n9742 & ~n9747;
  assign n9749 = ~n9741 & ~n9748;
  assign n9750 = ~n9740 & ~n9749;
  assign n9751 = ~n9739 & ~n9750;
  assign n9752 = ~n9738 & ~n9751;
  assign n9753 = ~n9737 & ~n9752;
  assign n9754 = ~n9736 & ~n9753;
  assign n9755 = ~n9735 & ~n9754;
  assign n9756 = ~n9734 & ~n9755;
  assign n9757 = ~pi184 & pi272;
  assign n9758 = pi183 & ~n9757;
  assign n9759 = ~n9756 & n9758;
  assign n9760 = pi271 & ~n9759;
  assign n9761 = ~n9756 & ~n9757;
  assign n9762 = ~pi183 & ~n9761;
  assign n9763 = ~n9760 & ~n9762;
  assign n9764 = pi184 & ~pi248;
  assign n9765 = ~pi185 & pi249;
  assign n9766 = pi185 & ~pi249;
  assign n9767 = ~pi186 & pi250;
  assign n9768 = pi186 & ~pi250;
  assign n9769 = ~pi187 & pi251;
  assign n9770 = pi187 & ~pi251;
  assign n9771 = ~pi188 & pi252;
  assign n9772 = pi188 & ~pi252;
  assign n9773 = pi190 & ~pi254;
  assign n9774 = pi189 & ~pi253;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = ~pi189 & pi253;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = ~n9772 & ~n9777;
  assign n9779 = ~n9771 & ~n9778;
  assign n9780 = ~n9770 & ~n9779;
  assign n9781 = ~n9769 & ~n9780;
  assign n9782 = ~n9768 & ~n9781;
  assign n9783 = ~n9767 & ~n9782;
  assign n9784 = ~n9766 & ~n9783;
  assign n9785 = ~n9765 & ~n9784;
  assign n9786 = ~n9764 & ~n9785;
  assign n9787 = ~pi184 & pi248;
  assign n9788 = pi183 & ~n9787;
  assign n9789 = ~n9786 & n9788;
  assign n9790 = pi247 & ~n9789;
  assign n9791 = ~n9786 & ~n9787;
  assign n9792 = ~pi183 & ~n9791;
  assign n9793 = ~n9790 & ~n9792;
  assign n9794 = ~n9763 & ~n9793;
  assign n9795 = pi184 & ~pi240;
  assign n9796 = ~pi185 & pi241;
  assign n9797 = pi185 & ~pi241;
  assign n9798 = ~pi186 & pi242;
  assign n9799 = pi186 & ~pi242;
  assign n9800 = ~pi187 & pi243;
  assign n9801 = pi187 & ~pi243;
  assign n9802 = ~pi188 & pi244;
  assign n9803 = pi188 & ~pi244;
  assign n9804 = pi190 & ~pi246;
  assign n9805 = pi189 & ~pi245;
  assign n9806 = ~n9804 & ~n9805;
  assign n9807 = ~pi189 & pi245;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = ~n9803 & ~n9808;
  assign n9810 = ~n9802 & ~n9809;
  assign n9811 = ~n9801 & ~n9810;
  assign n9812 = ~n9800 & ~n9811;
  assign n9813 = ~n9799 & ~n9812;
  assign n9814 = ~n9798 & ~n9813;
  assign n9815 = ~n9797 & ~n9814;
  assign n9816 = ~n9796 & ~n9815;
  assign n9817 = ~n9795 & ~n9816;
  assign n9818 = ~pi184 & pi240;
  assign n9819 = pi183 & ~n9818;
  assign n9820 = ~n9817 & n9819;
  assign n9821 = pi239 & ~n9820;
  assign n9822 = ~n9817 & ~n9818;
  assign n9823 = ~pi183 & ~n9822;
  assign n9824 = ~n9821 & ~n9823;
  assign n9825 = pi184 & ~pi256;
  assign n9826 = ~pi185 & pi257;
  assign n9827 = pi185 & ~pi257;
  assign n9828 = ~pi186 & pi258;
  assign n9829 = pi186 & ~pi258;
  assign n9830 = ~pi187 & pi259;
  assign n9831 = pi187 & ~pi259;
  assign n9832 = ~pi188 & pi260;
  assign n9833 = pi188 & ~pi260;
  assign n9834 = pi190 & ~pi262;
  assign n9835 = pi189 & ~pi261;
  assign n9836 = ~n9834 & ~n9835;
  assign n9837 = ~pi189 & pi261;
  assign n9838 = ~n9836 & ~n9837;
  assign n9839 = ~n9833 & ~n9838;
  assign n9840 = ~n9832 & ~n9839;
  assign n9841 = ~n9831 & ~n9840;
  assign n9842 = ~n9830 & ~n9841;
  assign n9843 = ~n9829 & ~n9842;
  assign n9844 = ~n9828 & ~n9843;
  assign n9845 = ~n9827 & ~n9844;
  assign n9846 = ~n9826 & ~n9845;
  assign n9847 = ~n9825 & ~n9846;
  assign n9848 = ~pi184 & pi256;
  assign n9849 = pi183 & ~n9848;
  assign n9850 = ~n9847 & n9849;
  assign n9851 = pi255 & ~n9850;
  assign n9852 = ~n9847 & ~n9848;
  assign n9853 = ~pi183 & ~n9852;
  assign n9854 = ~n9851 & ~n9853;
  assign n9855 = ~n9824 & ~n9854;
  assign n9856 = n9794 & n9855;
  assign n9857 = ~n7299 & ~n8705;
  assign n9858 = ~n8634 & n9857;
  assign n9859 = ~n6433 & ~n7240;
  assign n9860 = n6740 & n9859;
  assign n9861 = ~n4649 & ~n5499;
  assign n9862 = n5757 & n9861;
  assign n9863 = n9860 & n9862;
  assign n9864 = n9858 & n9863;
  assign n9865 = ~n1087 & ~n2052;
  assign n9866 = n3812 & n9865;
  assign n9867 = ~n1404 & ~n1620;
  assign n9868 = n5713 & n9867;
  assign n9869 = n9866 & n9868;
  assign n9870 = ~n3256 & ~n3496;
  assign n9871 = ~n2425 & ~n2694;
  assign n9872 = n9870 & n9871;
  assign n9873 = n3941 & n4849;
  assign n9874 = n9872 & n9873;
  assign n9875 = n9869 & n9874;
  assign n9876 = n3861 & n9875;
  assign n9877 = n9864 & n9876;
  assign n9878 = ~n1172 & n9877;
  assign n9879 = ~n1114 & n9878;
  assign n9880 = ~n996 & n9879;
  assign n9881 = ~n500 & n9880;
  assign n9882 = n2316 & n9881;
  assign n9883 = n7608 & n9882;
  assign n9884 = pi184 & ~pi264;
  assign n9885 = ~pi185 & pi265;
  assign n9886 = pi185 & ~pi265;
  assign n9887 = ~pi186 & pi266;
  assign n9888 = pi186 & ~pi266;
  assign n9889 = ~pi187 & pi267;
  assign n9890 = pi187 & ~pi267;
  assign n9891 = ~pi188 & pi268;
  assign n9892 = pi188 & ~pi268;
  assign n9893 = pi190 & ~pi270;
  assign n9894 = pi189 & ~pi269;
  assign n9895 = ~n9893 & ~n9894;
  assign n9896 = ~pi189 & pi269;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~n9892 & ~n9897;
  assign n9899 = ~n9891 & ~n9898;
  assign n9900 = ~n9890 & ~n9899;
  assign n9901 = ~n9889 & ~n9900;
  assign n9902 = ~n9888 & ~n9901;
  assign n9903 = ~n9887 & ~n9902;
  assign n9904 = ~n9886 & ~n9903;
  assign n9905 = ~n9885 & ~n9904;
  assign n9906 = ~n9884 & ~n9905;
  assign n9907 = ~pi184 & pi264;
  assign n9908 = pi183 & ~n9907;
  assign n9909 = ~n9906 & n9908;
  assign n9910 = pi263 & ~n9909;
  assign n9911 = ~n9906 & ~n9907;
  assign n9912 = ~pi183 & ~n9911;
  assign n9913 = ~n9910 & ~n9912;
  assign n9914 = ~n1648 & n4786;
  assign n9915 = ~n9913 & n9914;
  assign n9916 = n9883 & n9915;
  assign n9917 = n9856 & n9916;
  assign n9918 = n9733 & n9917;
  assign n9919 = ~n7236 & n9918;
  assign n9920 = ~n6137 & n9919;
  assign n9921 = n6193 & n9920;
  assign n9922 = n6134 & n9921;
  assign n9923 = ~n8867 & n9922;
  assign n9924 = ~n7235 & n9923;
  assign n9925 = n7296 & n9924;
  assign n9926 = n7231 & n9925;
  assign n9927 = ~n8866 & n9926;
  assign n9928 = n8898 & n9927;
  assign n9929 = n8863 & n9928;
  assign n9930 = ~n9533 & ~n9929;
  assign n9931 = n8733 & ~n8900;
  assign n9932 = ~n9300 & ~n9374;
  assign n9933 = ~n9931 & n9932;
  assign n9934 = ~n8603 & ~n8633;
  assign n9935 = ~n8455 & ~n8662;
  assign n9936 = n9934 & n9935;
  assign n9937 = ~n8762 & ~n8792;
  assign n9938 = ~n8574 & ~n8821;
  assign n9939 = n9937 & n9938;
  assign n9940 = n9936 & n9939;
  assign n9941 = ~n8484 & ~n8514;
  assign n9942 = ~n8543 & n9941;
  assign n9943 = ~n8426 & n9942;
  assign n9944 = n9940 & n9943;
  assign n9945 = ~n8834 & n9944;
  assign n9946 = ~n9185 & n9945;
  assign n9947 = ~n9207 & n9946;
  assign n9948 = ~n9458 & n9947;
  assign n9949 = ~n3679 & ~n3940;
  assign n9950 = ~n4001 & n9949;
  assign n9951 = ~n5043 & n9950;
  assign n9952 = ~n5943 & n9951;
  assign n9953 = ~n6951 & n9952;
  assign n9954 = ~n8037 & n9953;
  assign n9955 = ~n9515 & ~n9954;
  assign n9956 = n9948 & n9955;
  assign n9957 = n9933 & n9956;
  assign n9958 = ~n1026 & ~n1372;
  assign n9959 = ~n2243 & n9958;
  assign n9960 = ~n3104 & n9959;
  assign n9961 = ~n3971 & n9960;
  assign n9962 = ~n4872 & n9961;
  assign n9963 = ~n5801 & n9962;
  assign n9964 = ~n6739 & n9963;
  assign n9965 = ~n7807 & n9964;
  assign n9966 = ~n8989 & n9965;
  assign n9967 = ~n4370 & ~n4817;
  assign n9968 = ~n4902 & n9967;
  assign n9969 = ~n6001 & n9968;
  assign n9970 = ~n7014 & n9969;
  assign n9971 = ~n8114 & n9970;
  assign n9972 = ~n7534 & ~n7869;
  assign n9973 = ~n8346 & n9972;
  assign n9974 = ~n9971 & ~n9973;
  assign n9975 = ~n9966 & n9974;
  assign n9976 = ~n2842 & ~n3066;
  assign n9977 = ~n3983 & n9976;
  assign n9978 = ~n4024 & n9977;
  assign n9979 = ~n4999 & n9978;
  assign n9980 = ~n5827 & n9979;
  assign n9981 = ~n6893 & n9980;
  assign n9982 = ~n7890 & n9981;
  assign n9983 = ~n6432 & ~n6784;
  assign n9984 = ~n7158 & n9983;
  assign n9985 = ~n8250 & n9984;
  assign n9986 = ~n9982 & ~n9985;
  assign n9987 = ~n2020 & ~n2242;
  assign n9988 = ~n3095 & n9987;
  assign n9989 = ~n3997 & n9988;
  assign n9990 = ~n4837 & n9989;
  assign n9991 = ~n5822 & n9990;
  assign n9992 = ~n6820 & n9991;
  assign n9993 = ~n7785 & n9992;
  assign n9994 = ~n9027 & n9993;
  assign n9995 = ~n5259 & ~n5808;
  assign n9996 = ~n6056 & n9995;
  assign n9997 = ~n7073 & n9996;
  assign n9998 = ~n8179 & n9997;
  assign n9999 = ~n9994 & ~n9998;
  assign n10000 = n9986 & n9999;
  assign n10001 = n9975 & n10000;
  assign n10002 = n9957 & n10001;
  assign n10003 = ~n1897 & ~n2242;
  assign n10004 = ~n3095 & n10003;
  assign n10005 = ~n3997 & n10004;
  assign n10006 = ~n4837 & n10005;
  assign n10007 = ~n5822 & n10006;
  assign n10008 = ~n6820 & n10007;
  assign n10009 = ~n7785 & n10008;
  assign n10010 = ~n9027 & n10009;
  assign n10011 = ~n7595 & ~n7869;
  assign n10012 = ~n8346 & n10011;
  assign n10013 = ~n3024 & ~n3066;
  assign n10014 = ~n3983 & n10013;
  assign n10015 = ~n4024 & n10014;
  assign n10016 = ~n4999 & n10015;
  assign n10017 = ~n5827 & n10016;
  assign n10018 = ~n6893 & n10017;
  assign n10019 = ~n7890 & n10018;
  assign n10020 = ~n10012 & ~n10019;
  assign n10021 = ~n10010 & n10020;
  assign n10022 = ~n4192 & ~n4817;
  assign n10023 = ~n4902 & n10022;
  assign n10024 = ~n6001 & n10023;
  assign n10025 = ~n7014 & n10024;
  assign n10026 = ~n8114 & n10025;
  assign n10027 = ~n8426 & ~n8834;
  assign n10028 = n6677 & n7279;
  assign n10029 = n8879 & n10028;
  assign n10030 = n4786 & n9654;
  assign n10031 = n2316 & n8876;
  assign n10032 = n7608 & n10031;
  assign n10033 = n10030 & n10032;
  assign n10034 = n10029 & n10033;
  assign n10035 = ~n7236 & n10034;
  assign n10036 = ~n6137 & n10035;
  assign n10037 = n6193 & n10036;
  assign n10038 = n6134 & n10037;
  assign n10039 = ~n8867 & n10038;
  assign n10040 = ~n7235 & n10039;
  assign n10041 = n7296 & n10040;
  assign n10042 = n7231 & n10041;
  assign n10043 = ~n10027 & n10042;
  assign n10044 = ~n8866 & n10043;
  assign n10045 = n8898 & n10044;
  assign n10046 = n8863 & n10045;
  assign n10047 = ~n10026 & n10046;
  assign n10048 = ~n5170 & ~n5808;
  assign n10049 = ~n6056 & n10048;
  assign n10050 = ~n7073 & n10049;
  assign n10051 = ~n8179 & n10050;
  assign n10052 = ~n1270 & ~n1372;
  assign n10053 = ~n2243 & n10052;
  assign n10054 = ~n3104 & n10053;
  assign n10055 = ~n3971 & n10054;
  assign n10056 = ~n4872 & n10055;
  assign n10057 = ~n5801 & n10056;
  assign n10058 = ~n6739 & n10057;
  assign n10059 = ~n7807 & n10058;
  assign n10060 = ~n8989 & n10059;
  assign n10061 = ~n10051 & ~n10060;
  assign n10062 = ~n6224 & ~n6784;
  assign n10063 = ~n7158 & n10062;
  assign n10064 = ~n8250 & n10063;
  assign n10065 = ~n3464 & ~n3940;
  assign n10066 = ~n4001 & n10065;
  assign n10067 = ~n5043 & n10066;
  assign n10068 = ~n5943 & n10067;
  assign n10069 = ~n6951 & n10068;
  assign n10070 = ~n8037 & n10069;
  assign n10071 = ~n10064 & ~n10070;
  assign n10072 = n10061 & n10071;
  assign n10073 = n10047 & n10072;
  assign n10074 = n10021 & n10073;
  assign n10075 = ~n8179 & n8384;
  assign n10076 = ~n8114 & n8380;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = ~n8037 & n8381;
  assign n10079 = ~n7890 & n8385;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = n10077 & n10080;
  assign n10082 = n8388 & ~n8989;
  assign n10083 = n8387 & ~n9027;
  assign n10084 = ~n10082 & ~n10083;
  assign n10085 = ~n8250 & n8379;
  assign n10086 = ~n8346 & n8391;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = n10084 & n10087;
  assign n10089 = ~po161 & ~n9185;
  assign n10090 = ~n8397 & n10089;
  assign n10091 = ~n9458 & n10090;
  assign n10092 = n9443 & n10091;
  assign n10093 = n10088 & n10092;
  assign n10094 = n10081 & n10093;
  assign n10095 = ~n10074 & ~n10094;
  assign n10096 = ~n10002 & n10095;
  assign po169 = ~n9930 | ~n10096;
  assign n10098 = ~n9510 & ~po169;
  assign n10099 = pi020 & ~n501;
  assign n10100 = n5714 & n10099;
  assign n10101 = n5719 & n10100;
  assign n10102 = n8912 & n10101;
  assign n10103 = ~n1172 & n10102;
  assign n10104 = ~n996 & n10103;
  assign n10105 = ~n2306 & n10104;
  assign n10106 = ~n500 & n10105;
  assign n10107 = n2316 & n10106;
  assign n10108 = n7608 & n10107;
  assign n10109 = n10030 & n10108;
  assign n10110 = n10029 & n10109;
  assign n10111 = ~n7236 & n10110;
  assign n10112 = ~n6137 & n10111;
  assign n10113 = n6193 & n10112;
  assign n10114 = n6134 & n10113;
  assign n10115 = ~n8867 & n10114;
  assign n10116 = ~n7235 & n10115;
  assign n10117 = n7296 & n10116;
  assign n10118 = n7231 & n10117;
  assign n10119 = ~n10027 & n10118;
  assign n10120 = ~n8866 & n10119;
  assign n10121 = n8898 & n10120;
  assign n10122 = n8863 & n10121;
  assign n10123 = ~n10026 & n10122;
  assign n10124 = n10072 & n10123;
  assign n10125 = n10021 & n10124;
  assign n10126 = ~n6433 & ~n7299;
  assign n10127 = ~n8634 & ~n8705;
  assign n10128 = n10126 & n10127;
  assign n10129 = n4796 & n9861;
  assign n10130 = n7242 & n10129;
  assign n10131 = n10128 & n10130;
  assign n10132 = pi019 & ~n501;
  assign n10133 = n9865 & n9867;
  assign n10134 = n10132 & n10133;
  assign n10135 = n4790 & n8941;
  assign n10136 = n3810 & n4795;
  assign n10137 = n9872 & n10136;
  assign n10138 = n10135 & n10137;
  assign n10139 = n10134 & n10138;
  assign n10140 = n10131 & n10139;
  assign n10141 = ~n1172 & n10140;
  assign n10142 = ~n1114 & n10141;
  assign n10143 = ~n996 & n10142;
  assign n10144 = ~n500 & n10143;
  assign n10145 = n2316 & n10144;
  assign n10146 = n7608 & n10145;
  assign n10147 = n9915 & n10146;
  assign n10148 = n9856 & n10147;
  assign n10149 = n9733 & n10148;
  assign n10150 = ~n7236 & n10149;
  assign n10151 = ~n6137 & n10150;
  assign n10152 = n6193 & n10151;
  assign n10153 = n6134 & n10152;
  assign n10154 = ~n8867 & n10153;
  assign n10155 = ~n7235 & n10154;
  assign n10156 = n7296 & n10155;
  assign n10157 = n7231 & n10156;
  assign n10158 = ~n8866 & n10157;
  assign n10159 = n8898 & n10158;
  assign n10160 = n8863 & n10159;
  assign n10161 = ~n10125 & ~n10160;
  assign n10162 = pi016 & ~po161;
  assign n10163 = ~n9185 & n10162;
  assign n10164 = ~n8397 & n10163;
  assign n10165 = ~n9458 & n10164;
  assign n10166 = n9443 & n10165;
  assign n10167 = n10088 & n10166;
  assign n10168 = n10081 & n10167;
  assign n10169 = pi017 & ~n8762;
  assign n10170 = n8822 & n10169;
  assign n10171 = n8664 & n10170;
  assign n10172 = ~n8426 & n8545;
  assign n10173 = n10171 & n10172;
  assign n10174 = ~n8834 & n10173;
  assign n10175 = ~n9185 & n10174;
  assign n10176 = ~n9207 & n10175;
  assign n10177 = ~n9458 & n10176;
  assign n10178 = n9955 & n10177;
  assign n10179 = n9933 & n10178;
  assign n10180 = n10001 & n10179;
  assign n10181 = pi018 & ~n9511;
  assign n10182 = ~n8900 & n10181;
  assign n10183 = ~n9185 & n10182;
  assign n10184 = ~n9458 & n10183;
  assign n10185 = n9517 & n10184;
  assign n10186 = n9443 & n10185;
  assign n10187 = n9532 & n10186;
  assign n10188 = ~n10180 & ~n10187;
  assign n10189 = ~n10168 & n10188;
  assign n10190 = n10161 & n10189;
  assign po010 = n10098 | ~n10190;
  assign n10192 = n9102 & ~n9414;
  assign n10193 = n9112 & ~n9485;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = n3024 & ~n10074;
  assign n10196 = n9099 & ~n9200;
  assign n10197 = ~n10195 & ~n10196;
  assign n10198 = n10194 & n10197;
  assign n10199 = n9105 & ~n9215;
  assign n10200 = n9106 & ~n9381;
  assign n10201 = n9109 & ~n9307;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = ~n10199 & n10202;
  assign n10204 = n9101 & ~n9344;
  assign n10205 = n9113 & ~n9160;
  assign n10206 = n2453 & ~n9929;
  assign n10207 = ~n2424 & ~n2483;
  assign n10208 = n2632 & n10207;
  assign n10209 = n2573 & n10208;
  assign n10210 = n9137 & n10209;
  assign n10211 = ~n3066 & n10210;
  assign n10212 = ~n3983 & n10211;
  assign n10213 = ~n4003 & n10212;
  assign n10214 = ~n4024 & n10213;
  assign n10215 = ~n4999 & n10214;
  assign n10216 = ~n5827 & n10215;
  assign n10217 = ~n6893 & n10216;
  assign n10218 = ~n7890 & n10217;
  assign n10219 = ~n10206 & n10218;
  assign n10220 = ~n10205 & n10219;
  assign n10221 = ~n9131 & n10220;
  assign n10222 = ~n10204 & n10221;
  assign n10223 = n10203 & n10222;
  assign n10224 = n10198 & n10223;
  assign n10225 = n9114 & ~n10002;
  assign n10226 = ~n1649 & ~n2206;
  assign n10227 = n3088 & n10226;
  assign n10228 = ~n1897 & n10227;
  assign n10229 = n4955 & n7909;
  assign n10230 = n10228 & n10229;
  assign n10231 = ~n2242 & n10230;
  assign n10232 = ~n3095 & n10231;
  assign n10233 = ~n3997 & n10232;
  assign n10234 = ~n4003 & n10233;
  assign n10235 = ~n4837 & n10234;
  assign n10236 = ~n5822 & n10235;
  assign n10237 = ~n6820 & n10236;
  assign n10238 = ~n7785 & n10237;
  assign n10239 = ~n9029 & n10238;
  assign n10240 = ~n9028 & n10239;
  assign n10241 = ~n9027 & n10240;
  assign n10242 = ~n9010 & n10241;
  assign n10243 = n9009 & n10242;
  assign n10244 = n9002 & n10243;
  assign n10245 = n8995 & n10244;
  assign n10246 = n9094 & ~n10245;
  assign n10247 = n9095 & ~n9453;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = ~n10225 & n10248;
  assign n10250 = n9108 & ~n9533;
  assign n10251 = n9098 & ~n9276;
  assign n10252 = ~n10250 & ~n10251;
  assign n10253 = n9091 & ~n10094;
  assign n10254 = ~n1115 & ~n1208;
  assign n10255 = n4920 & n10254;
  assign n10256 = ~n1270 & n10255;
  assign n10257 = n4932 & n10256;
  assign n10258 = ~n1372 & n10257;
  assign n10259 = ~n2243 & n10258;
  assign n10260 = ~n3104 & n10259;
  assign n10261 = ~n3837 & n10260;
  assign n10262 = ~n3971 & n10261;
  assign n10263 = ~n4872 & n10262;
  assign n10264 = ~n5801 & n10263;
  assign n10265 = ~n6739 & n10264;
  assign n10266 = ~n7807 & n10265;
  assign n10267 = ~n9070 & n10266;
  assign n10268 = ~n9069 & n10267;
  assign n10269 = ~n9068 & n10268;
  assign n10270 = ~n9067 & n10269;
  assign n10271 = n9066 & n10270;
  assign n10272 = n9060 & n10271;
  assign n10273 = n9053 & n10272;
  assign n10274 = n9092 & ~n10273;
  assign n10275 = ~n10253 & ~n10274;
  assign n10276 = n10252 & n10275;
  assign n10277 = n10249 & n10276;
  assign n10278 = n10224 & n10277;
  assign n10279 = n9048 & ~n9131;
  assign n10280 = n9058 & ~n9344;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n9047 & ~n9200;
  assign n10283 = n9062 & ~n9533;
  assign n10284 = ~n10282 & ~n10283;
  assign n10285 = n10281 & n10284;
  assign n10286 = n9068 & ~n9215;
  assign n10287 = n9061 & ~n9381;
  assign n10288 = n9064 & ~n9307;
  assign n10289 = ~n10287 & ~n10288;
  assign n10290 = ~n10286 & n10289;
  assign n10291 = n1270 & ~n10074;
  assign n10292 = n9069 & ~n9160;
  assign n10293 = n1115 & ~n9929;
  assign n10294 = pi001 & ~n1208;
  assign n10295 = n4920 & n10294;
  assign n10296 = n4931 & n10295;
  assign n10297 = n4928 & n10296;
  assign n10298 = ~n1372 & n10297;
  assign n10299 = ~n2243 & n10298;
  assign n10300 = ~n3104 & n10299;
  assign n10301 = ~n3971 & n10300;
  assign n10302 = ~n4003 & n10301;
  assign n10303 = ~n4872 & n10302;
  assign n10304 = ~n5801 & n10303;
  assign n10305 = ~n6739 & n10304;
  assign n10306 = ~n7807 & n10305;
  assign n10307 = ~n8989 & n10306;
  assign n10308 = ~n10293 & n10307;
  assign n10309 = ~n10292 & n10308;
  assign n10310 = ~n10273 & n10309;
  assign n10311 = ~n10291 & n10310;
  assign n10312 = n10290 & n10311;
  assign n10313 = n10285 & n10312;
  assign n10314 = n9070 & ~n10002;
  assign n10315 = n9067 & ~n9485;
  assign n10316 = n9051 & ~n9453;
  assign n10317 = ~n10315 & ~n10316;
  assign n10318 = ~n10314 & n10317;
  assign n10319 = n9057 & ~n9414;
  assign n10320 = n9050 & ~n9276;
  assign n10321 = ~n10319 & ~n10320;
  assign n10322 = n9054 & ~n10094;
  assign n10323 = n9055 & ~n10245;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = n10321 & n10324;
  assign n10326 = n10318 & n10325;
  assign n10327 = n10313 & n10326;
  assign n10328 = n8997 & ~n9131;
  assign n10329 = n9010 & ~n9344;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = n8996 & ~n9200;
  assign n10332 = n9006 & ~n9533;
  assign n10333 = ~n10331 & ~n10332;
  assign n10334 = n10330 & n10333;
  assign n10335 = n9003 & ~n9215;
  assign n10336 = n9004 & ~n9381;
  assign n10337 = n9007 & ~n9307;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = ~n10335 & n10338;
  assign n10340 = n1897 & ~n10074;
  assign n10341 = n9028 & ~n9160;
  assign n10342 = n1649 & ~n9929;
  assign n10343 = n2255 & n4955;
  assign n10344 = n7909 & n10343;
  assign n10345 = ~n2242 & n10344;
  assign n10346 = ~n3095 & n10345;
  assign n10347 = ~n3997 & n10346;
  assign n10348 = ~n4003 & n10347;
  assign n10349 = ~n4837 & n10348;
  assign n10350 = ~n5822 & n10349;
  assign n10351 = ~n6820 & n10350;
  assign n10352 = ~n7785 & n10351;
  assign n10353 = ~n9027 & n10352;
  assign n10354 = ~n10342 & n10353;
  assign n10355 = ~n10341 & n10354;
  assign n10356 = ~n10245 & n10355;
  assign n10357 = ~n10340 & n10356;
  assign n10358 = n10339 & n10357;
  assign n10359 = n10334 & n10358;
  assign n10360 = n9029 & ~n10002;
  assign n10361 = n9000 & ~n9485;
  assign n10362 = n8993 & ~n9453;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = ~n10360 & n10363;
  assign n10365 = n8992 & ~n9414;
  assign n10366 = n8999 & ~n9276;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = n8968 & ~n10094;
  assign n10369 = n8990 & ~n10273;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = n10367 & n10370;
  assign n10372 = n10364 & n10371;
  assign n10373 = n10359 & n10372;
  assign n10374 = ~n10327 & ~n10373;
  assign n10375 = ~n10278 & n10374;
  assign n10376 = n2513 & n3852;
  assign n10377 = n9134 & n10376;
  assign n10378 = n9115 & n10377;
  assign n10379 = ~n3066 & n10378;
  assign n10380 = ~n3983 & n10379;
  assign n10381 = ~n4003 & n10380;
  assign n10382 = ~n4024 & n10381;
  assign n10383 = ~n4999 & n10382;
  assign n10384 = ~n5827 & n10383;
  assign n10385 = ~n6893 & n10384;
  assign n10386 = ~n7890 & n10385;
  assign n10387 = ~n10206 & n10386;
  assign n10388 = ~n10205 & n10387;
  assign n10389 = ~n9131 & n10388;
  assign n10390 = ~n10204 & n10389;
  assign n10391 = n10203 & n10390;
  assign n10392 = n10198 & n10391;
  assign n10393 = n10277 & n10392;
  assign n10394 = ~n9131 & n9154;
  assign n10395 = n9155 & ~n9160;
  assign n10396 = ~n10394 & n10395;
  assign n10397 = n9157 & ~n10245;
  assign n10398 = n9158 & ~n10273;
  assign n10399 = ~n10397 & ~n10398;
  assign n10400 = n10396 & n10399;
  assign n10401 = ~n10393 & ~n10400;
  assign n10402 = ~n10375 & n10401;
  assign n10403 = n9180 & ~n9533;
  assign n10404 = n9173 & ~n9344;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = n3464 & ~n10074;
  assign n10407 = ~n9131 & n9171;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = n10405 & n10408;
  assign n10410 = n9177 & ~n9215;
  assign n10411 = n9178 & ~n9381;
  assign n10412 = n9181 & ~n9307;
  assign n10413 = ~n10411 & ~n10412;
  assign n10414 = ~n10410 & n10413;
  assign n10415 = n9184 & ~n9414;
  assign n10416 = ~n9160 & n9185;
  assign n10417 = n3524 & ~n9929;
  assign n10418 = n3740 & n3951;
  assign n10419 = n9219 & n10418;
  assign n10420 = ~n3940 & n10419;
  assign n10421 = ~n4001 & n10420;
  assign n10422 = ~n5043 & n10421;
  assign n10423 = ~n5943 & n10422;
  assign n10424 = ~n6951 & n10423;
  assign n10425 = ~n8037 & n10424;
  assign n10426 = ~n10417 & n10425;
  assign n10427 = ~n10416 & n10426;
  assign n10428 = ~n9200 & n10427;
  assign n10429 = ~n10415 & n10428;
  assign n10430 = n10414 & n10429;
  assign n10431 = n10409 & n10430;
  assign n10432 = n9186 & ~n10002;
  assign n10433 = n9174 & ~n10245;
  assign n10434 = n9167 & ~n9453;
  assign n10435 = ~n10433 & ~n10434;
  assign n10436 = ~n10432 & n10435;
  assign n10437 = n9166 & ~n9485;
  assign n10438 = n9170 & ~n9276;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = n9164 & ~n10273;
  assign n10441 = n9163 & ~n10094;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = n10439 & n10442;
  assign n10444 = n10436 & n10443;
  assign n10445 = n10431 & n10444;
  assign n10446 = ~n9160 & n9201;
  assign n10447 = ~n10394 & n10446;
  assign n10448 = n10399 & n10447;
  assign n10449 = ~n10445 & ~n10448;
  assign n10450 = ~n10402 & n10449;
  assign n10451 = n9206 & ~n10273;
  assign n10452 = n9207 & ~n9215;
  assign n10453 = ~n10416 & n10452;
  assign n10454 = ~n10451 & n10453;
  assign n10455 = ~n9200 & n9210;
  assign n10456 = ~n9131 & n9211;
  assign n10457 = n9212 & ~n10245;
  assign n10458 = ~n10456 & ~n10457;
  assign n10459 = ~n10455 & n10458;
  assign n10460 = n10454 & n10459;
  assign n10461 = ~pi007 & ~n3710;
  assign n10462 = n4096 & n10461;
  assign n10463 = n4104 & n10462;
  assign n10464 = n8056 & n10463;
  assign n10465 = ~n3940 & n10464;
  assign n10466 = ~n4001 & n10465;
  assign n10467 = ~n5043 & n10466;
  assign n10468 = ~n5943 & n10467;
  assign n10469 = ~n6951 & n10468;
  assign n10470 = ~n8037 & n10469;
  assign n10471 = ~n10417 & n10470;
  assign n10472 = ~n10416 & n10471;
  assign n10473 = ~n9200 & n10472;
  assign n10474 = ~n10415 & n10473;
  assign n10475 = n10414 & n10474;
  assign n10476 = n10409 & n10475;
  assign n10477 = n10444 & n10476;
  assign n10478 = ~n10460 & ~n10477;
  assign n10479 = ~n10450 & n10478;
  assign n10480 = ~n9215 & n9236;
  assign n10481 = ~n10416 & n10480;
  assign n10482 = ~n10451 & n10481;
  assign n10483 = n10459 & n10482;
  assign n10484 = n9256 & ~n9533;
  assign n10485 = n9251 & ~n9414;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = n4192 & ~n10074;
  assign n10488 = ~n9131 & n9241;
  assign n10489 = ~n10487 & ~n10488;
  assign n10490 = n10486 & n10489;
  assign n10491 = n9257 & ~n9307;
  assign n10492 = n9254 & ~n9381;
  assign n10493 = ~n10452 & ~n10492;
  assign n10494 = ~n10491 & n10493;
  assign n10495 = ~n9200 & n9240;
  assign n10496 = n4677 & ~n9929;
  assign n10497 = n4491 & n4737;
  assign n10498 = n9281 & n10497;
  assign n10499 = ~n4817 & n10498;
  assign n10500 = ~n4902 & n10499;
  assign n10501 = ~n6001 & n10500;
  assign n10502 = ~n7014 & n10501;
  assign n10503 = ~n8114 & n10502;
  assign n10504 = ~n10496 & n10503;
  assign n10505 = ~n10416 & n10504;
  assign n10506 = ~n9276 & n10505;
  assign n10507 = ~n10495 & n10506;
  assign n10508 = n10494 & n10507;
  assign n10509 = n10490 & n10508;
  assign n10510 = n9261 & ~n10002;
  assign n10511 = n9260 & ~n10245;
  assign n10512 = n9247 & ~n10094;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = ~n10510 & n10513;
  assign n10515 = n9250 & ~n9485;
  assign n10516 = n9243 & ~n9344;
  assign n10517 = ~n10515 & ~n10516;
  assign n10518 = n9244 & ~n9453;
  assign n10519 = n9248 & ~n10273;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = n10517 & n10520;
  assign n10522 = n10514 & n10521;
  assign n10523 = n10509 & n10522;
  assign n10524 = ~n10483 & ~n10523;
  assign n10525 = ~n10479 & n10524;
  assign n10526 = ~pi009 & ~n4707;
  assign n10527 = n5083 & n10526;
  assign n10528 = n8096 & n10527;
  assign n10529 = n9263 & n10528;
  assign n10530 = ~n4817 & n10529;
  assign n10531 = ~n4902 & n10530;
  assign n10532 = ~n6001 & n10531;
  assign n10533 = ~n7014 & n10532;
  assign n10534 = ~n8114 & n10533;
  assign n10535 = ~n10496 & n10534;
  assign n10536 = ~n10416 & n10535;
  assign n10537 = ~n9276 & n10536;
  assign n10538 = ~n10495 & n10537;
  assign n10539 = n10494 & n10538;
  assign n10540 = n10490 & n10539;
  assign n10541 = n10522 & n10540;
  assign n10542 = n9295 & ~n10273;
  assign n10543 = ~n9131 & n9296;
  assign n10544 = n9297 & ~n10245;
  assign n10545 = ~n10543 & ~n10544;
  assign n10546 = ~n10542 & n10545;
  assign n10547 = n9300 & ~n9307;
  assign n10548 = ~n10416 & n10547;
  assign n10549 = ~n10452 & n10548;
  assign n10550 = ~n9200 & n9303;
  assign n10551 = ~n9276 & n9304;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = n10549 & n10552;
  assign n10554 = n10546 & n10553;
  assign n10555 = ~n10541 & ~n10554;
  assign n10556 = ~n10525 & n10555;
  assign n10557 = n9326 & ~n9533;
  assign n10558 = n9321 & ~n9414;
  assign n10559 = ~n10557 & ~n10558;
  assign n10560 = n5170 & ~n10074;
  assign n10561 = ~n9131 & n9311;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = n10559 & n10562;
  assign n10564 = ~n10452 & ~n10547;
  assign n10565 = n9325 & ~n9381;
  assign n10566 = n10564 & ~n10565;
  assign n10567 = ~n9200 & n9310;
  assign n10568 = n5527 & ~n9929;
  assign n10569 = n5438 & n9331;
  assign n10570 = n6040 & n10569;
  assign n10571 = ~n5808 & n10570;
  assign n10572 = ~n6056 & n10571;
  assign n10573 = ~n7073 & n10572;
  assign n10574 = ~n8179 & n10573;
  assign n10575 = ~n10568 & n10574;
  assign n10576 = ~n10416 & n10575;
  assign n10577 = ~n9344 & n10576;
  assign n10578 = ~n10567 & n10577;
  assign n10579 = n10566 & n10578;
  assign n10580 = n10563 & n10579;
  assign n10581 = n9330 & ~n10002;
  assign n10582 = n9329 & ~n10245;
  assign n10583 = n9317 & ~n10094;
  assign n10584 = ~n10582 & ~n10583;
  assign n10585 = ~n10581 & n10584;
  assign n10586 = n9320 & ~n9485;
  assign n10587 = ~n9276 & n9313;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = n9314 & ~n9453;
  assign n10590 = n9318 & ~n10273;
  assign n10591 = ~n10589 & ~n10590;
  assign n10592 = n10588 & n10591;
  assign n10593 = n10585 & n10592;
  assign n10594 = n10580 & n10593;
  assign n10595 = ~n9307 & n9345;
  assign n10596 = ~n10416 & n10595;
  assign n10597 = ~n10452 & n10596;
  assign n10598 = n10552 & n10597;
  assign n10599 = n10546 & n10598;
  assign n10600 = ~n10594 & ~n10599;
  assign n10601 = ~n10556 & n10600;
  assign n10602 = ~n5289 & n6073;
  assign n10603 = n9353 & n10602;
  assign n10604 = ~n5808 & n10603;
  assign n10605 = ~n6056 & n10604;
  assign n10606 = ~n7073 & n10605;
  assign n10607 = ~n8179 & n10606;
  assign n10608 = ~n10568 & n10607;
  assign n10609 = ~n10416 & n10608;
  assign n10610 = ~n9344 & n10609;
  assign n10611 = ~n10567 & n10610;
  assign n10612 = n10566 & n10611;
  assign n10613 = n10563 & n10612;
  assign n10614 = n10593 & n10613;
  assign n10615 = ~n9131 & n9367;
  assign n10616 = ~n9276 & n9368;
  assign n10617 = ~n10615 & ~n10616;
  assign n10618 = n9370 & ~n10273;
  assign n10619 = n9371 & ~n10245;
  assign n10620 = ~n10618 & ~n10619;
  assign n10621 = n10617 & n10620;
  assign n10622 = n9374 & ~n9381;
  assign n10623 = ~n10416 & n10622;
  assign n10624 = n10564 & n10623;
  assign n10625 = ~n9344 & n9377;
  assign n10626 = ~n9200 & n9378;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = n10624 & n10627;
  assign n10629 = n10621 & n10628;
  assign n10630 = ~n10614 & ~n10629;
  assign n10631 = ~n10601 & n10630;
  assign n10632 = ~n9344 & n9395;
  assign n10633 = n9398 & ~n9533;
  assign n10634 = ~n10632 & ~n10633;
  assign n10635 = n6224 & ~n10074;
  assign n10636 = ~n9131 & n9385;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 = n10634 & n10637;
  assign n10639 = ~n10452 & ~n10622;
  assign n10640 = ~n10547 & n10639;
  assign n10641 = ~n9276 & n9387;
  assign n10642 = n6461 & ~n9929;
  assign n10643 = n6343 & n8233;
  assign n10644 = n8236 & n10643;
  assign n10645 = ~n6784 & n10644;
  assign n10646 = ~n7158 & n10645;
  assign n10647 = ~n8250 & n10646;
  assign n10648 = ~n10642 & n10647;
  assign n10649 = ~n10416 & n10648;
  assign n10650 = ~n9414 & n10649;
  assign n10651 = ~n10641 & n10650;
  assign n10652 = n10640 & n10651;
  assign n10653 = n10638 & n10652;
  assign n10654 = n9402 & ~n10002;
  assign n10655 = n9401 & ~n10245;
  assign n10656 = n9391 & ~n10094;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10654 & n10657;
  assign n10659 = n9394 & ~n9485;
  assign n10660 = ~n9200 & n9384;
  assign n10661 = ~n10659 & ~n10660;
  assign n10662 = n9388 & ~n9453;
  assign n10663 = n9392 & ~n10273;
  assign n10664 = ~n10662 & ~n10663;
  assign n10665 = n10661 & n10664;
  assign n10666 = n10658 & n10665;
  assign n10667 = n10653 & n10666;
  assign n10668 = ~n9381 & n9415;
  assign n10669 = ~n10416 & n10668;
  assign n10670 = n10564 & n10669;
  assign n10671 = n10627 & n10670;
  assign n10672 = n10621 & n10671;
  assign n10673 = ~n10667 & ~n10672;
  assign n10674 = ~n10631 & n10673;
  assign n10675 = ~pi013 & ~n6313;
  assign n10676 = n7169 & n10675;
  assign n10677 = n7177 & n10676;
  assign n10678 = n8261 & n10677;
  assign n10679 = ~n6784 & n10678;
  assign n10680 = ~n7158 & n10679;
  assign n10681 = ~n8250 & n10680;
  assign n10682 = ~n10642 & n10681;
  assign n10683 = ~n10416 & n10682;
  assign n10684 = ~n9414 & n10683;
  assign n10685 = ~n10641 & n10684;
  assign n10686 = n10640 & n10685;
  assign n10687 = n10638 & n10686;
  assign n10688 = n10666 & n10687;
  assign n10689 = ~n9414 & n9436;
  assign n10690 = ~n9344 & n9437;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n9131 & n9439;
  assign n10693 = ~n9276 & n9440;
  assign n10694 = ~n10692 & ~n10693;
  assign n10695 = n10691 & n10694;
  assign n10696 = n9444 & ~n10273;
  assign n10697 = n9458 & ~n10416;
  assign n10698 = ~n9453 & n10697;
  assign n10699 = ~n10696 & n10698;
  assign n10700 = n9448 & ~n10245;
  assign n10701 = ~n9200 & n9449;
  assign n10702 = ~n10700 & ~n10701;
  assign n10703 = n10699 & n10702;
  assign n10704 = n10640 & n10703;
  assign n10705 = n10695 & n10704;
  assign n10706 = ~n9200 & n9454;
  assign n10707 = ~n9276 & n9457;
  assign n10708 = ~n10706 & ~n10707;
  assign n10709 = ~n9344 & n9465;
  assign n10710 = n7595 & ~n10074;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = n10708 & n10711;
  assign n10713 = ~n9453 & n9458;
  assign n10714 = n7327 & ~n9929;
  assign n10715 = ~n7356 & ~n7505;
  assign n10716 = n7416 & n10715;
  assign n10717 = n7476 & n7752;
  assign n10718 = n7693 & n10717;
  assign n10719 = n10716 & n10718;
  assign n10720 = ~n7869 & n10719;
  assign n10721 = ~n8346 & n10720;
  assign n10722 = ~n10714 & n10721;
  assign n10723 = ~n10416 & n10722;
  assign n10724 = ~n9485 & n10723;
  assign n10725 = ~n10713 & n10724;
  assign n10726 = n10640 & n10725;
  assign n10727 = n10712 & n10726;
  assign n10728 = n9472 & ~n10002;
  assign n10729 = ~n9414 & n9464;
  assign n10730 = n9462 & ~n10273;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = ~n10728 & n10731;
  assign n10733 = n9468 & ~n9533;
  assign n10734 = ~n9131 & n9455;
  assign n10735 = ~n10733 & ~n10734;
  assign n10736 = n9461 & ~n10094;
  assign n10737 = n9471 & ~n10245;
  assign n10738 = ~n10736 & ~n10737;
  assign n10739 = n10735 & n10738;
  assign n10740 = n10732 & n10739;
  assign n10741 = n10727 & n10740;
  assign n10742 = ~n10705 & ~n10741;
  assign n10743 = ~n10688 & n10742;
  assign n10744 = ~n10674 & n10743;
  assign n10745 = ~n8291 & n9489;
  assign n10746 = ~n10416 & n10745;
  assign n10747 = ~n9453 & n10746;
  assign n10748 = ~n10696 & n10747;
  assign n10749 = n10702 & n10748;
  assign n10750 = n10640 & n10749;
  assign n10751 = n10695 & n10750;
  assign n10752 = n8363 & n9498;
  assign n10753 = ~n7869 & n10752;
  assign n10754 = ~n8346 & n10753;
  assign n10755 = ~n10714 & n10754;
  assign n10756 = ~n10416 & n10755;
  assign n10757 = ~n9485 & n10756;
  assign n10758 = ~n10713 & n10757;
  assign n10759 = n10640 & n10758;
  assign n10760 = n10712 & n10759;
  assign n10761 = n10740 & n10760;
  assign n10762 = ~n10751 & ~n10761;
  assign n10763 = ~n10744 & n10762;
  assign n10764 = ~n9344 & n9521;
  assign n10765 = ~n8900 & ~n10416;
  assign n10766 = ~n9533 & n10765;
  assign n10767 = ~n10764 & n10766;
  assign n10768 = ~n9414 & n9528;
  assign n10769 = ~n9485 & n9525;
  assign n10770 = ~n10768 & ~n10769;
  assign n10771 = n10767 & n10770;
  assign n10772 = n10640 & n10771;
  assign n10773 = ~n9276 & n9520;
  assign n10774 = ~n10713 & ~n10773;
  assign n10775 = n9516 & ~n10245;
  assign n10776 = ~n9131 & n9529;
  assign n10777 = ~n10775 & ~n10776;
  assign n10778 = n10774 & n10777;
  assign n10779 = n9511 & ~n10002;
  assign n10780 = n9515 & ~n10094;
  assign n10781 = ~n10779 & ~n10780;
  assign n10782 = n9526 & ~n10273;
  assign n10783 = ~n9200 & n9522;
  assign n10784 = ~n10782 & ~n10783;
  assign n10785 = n10781 & n10784;
  assign n10786 = n10778 & n10785;
  assign n10787 = n10772 & n10786;
  assign n10788 = ~n9562 & ~n9929;
  assign n10789 = pi200 & ~pi208;
  assign n10790 = ~pi201 & pi209;
  assign n10791 = pi201 & ~pi209;
  assign n10792 = ~pi202 & pi210;
  assign n10793 = pi202 & ~pi210;
  assign n10794 = ~pi203 & pi211;
  assign n10795 = pi203 & ~pi211;
  assign n10796 = ~pi205 & pi213;
  assign n10797 = pi206 & ~pi214;
  assign n10798 = ~n10796 & n10797;
  assign n10799 = pi205 & ~pi213;
  assign n10800 = pi204 & ~pi212;
  assign n10801 = ~n10799 & ~n10800;
  assign n10802 = ~n10798 & n10801;
  assign n10803 = ~pi204 & pi212;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = ~n10795 & ~n10804;
  assign n10806 = ~n10794 & ~n10805;
  assign n10807 = ~n10793 & ~n10806;
  assign n10808 = ~n10792 & ~n10807;
  assign n10809 = ~n10791 & ~n10808;
  assign n10810 = ~n10790 & ~n10809;
  assign n10811 = ~n10789 & ~n10810;
  assign n10812 = ~pi200 & pi208;
  assign n10813 = pi199 & ~n10812;
  assign n10814 = ~n10811 & n10813;
  assign n10815 = pi207 & ~n10814;
  assign n10816 = ~n10811 & ~n10812;
  assign n10817 = ~pi199 & ~n10816;
  assign n10818 = ~n10815 & ~n10817;
  assign n10819 = n9654 & n10818;
  assign n10820 = ~n2080 & ~n2142;
  assign n10821 = n3822 & n10820;
  assign n10822 = n4787 & n10821;
  assign n10823 = n10819 & n10822;
  assign n10824 = ~n7414 & ~n8732;
  assign n10825 = ~n8791 & n10824;
  assign n10826 = ~n6341 & ~n7277;
  assign n10827 = n6181 & n10826;
  assign n10828 = ~n4607 & ~n5288;
  assign n10829 = n5732 & n10828;
  assign n10830 = n10827 & n10829;
  assign n10831 = n10825 & n10830;
  assign n10832 = ~n7387 & ~n8705;
  assign n10833 = ~n8764 & n10832;
  assign n10834 = ~n6314 & ~n7240;
  assign n10835 = n6740 & n10834;
  assign n10836 = ~n4580 & ~n5261;
  assign n10837 = n5757 & n10836;
  assign n10838 = n10835 & n10837;
  assign n10839 = n10833 & n10838;
  assign n10840 = ~n628 & ~n969;
  assign n10841 = ~n1145 & ~n2114;
  assign n10842 = n10840 & n10841;
  assign n10843 = n5718 & n10842;
  assign n10844 = ~n3256 & ~n3345;
  assign n10845 = ~n2484 & ~n2694;
  assign n10846 = n10844 & n10845;
  assign n10847 = n9873 & n10846;
  assign n10848 = n10843 & n10847;
  assign n10849 = n3861 & n10848;
  assign n10850 = n10839 & n10849;
  assign n10851 = ~n1172 & n10850;
  assign n10852 = ~n996 & n10851;
  assign n10853 = ~n2306 & n10852;
  assign n10854 = ~n500 & n10853;
  assign n10855 = ~n532 & ~n656;
  assign n10856 = n10854 & n10855;
  assign n10857 = ~n3283 & ~n3372;
  assign n10858 = ~n2511 & ~n2721;
  assign n10859 = n10857 & n10858;
  assign n10860 = n7601 & n10859;
  assign n10861 = n10856 & n10860;
  assign n10862 = n10831 & n10861;
  assign n10863 = n10823 & n10862;
  assign n10864 = ~n7236 & n10863;
  assign n10865 = ~n6137 & n10864;
  assign n10866 = n6193 & n10865;
  assign n10867 = n6134 & n10866;
  assign n10868 = ~n8867 & n10867;
  assign n10869 = ~n7235 & n10868;
  assign n10870 = n7296 & n10869;
  assign n10871 = n7231 & n10870;
  assign n10872 = ~n10027 & n10871;
  assign n10873 = ~n8866 & n10872;
  assign n10874 = n8898 & n10873;
  assign n10875 = n8863 & n10874;
  assign n10876 = ~n10788 & n10875;
  assign n10877 = ~n10026 & n10876;
  assign n10878 = n10072 & n10877;
  assign n10879 = n10021 & n10878;
  assign n10880 = pi200 & ~pi232;
  assign n10881 = ~pi201 & pi233;
  assign n10882 = pi201 & ~pi233;
  assign n10883 = ~pi202 & pi234;
  assign n10884 = pi202 & ~pi234;
  assign n10885 = ~pi203 & pi235;
  assign n10886 = pi203 & ~pi235;
  assign n10887 = ~pi205 & pi237;
  assign n10888 = pi206 & ~pi238;
  assign n10889 = ~n10887 & n10888;
  assign n10890 = pi205 & ~pi237;
  assign n10891 = pi204 & ~pi236;
  assign n10892 = ~n10890 & ~n10891;
  assign n10893 = ~n10889 & n10892;
  assign n10894 = ~pi204 & pi236;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = ~n10886 & ~n10895;
  assign n10897 = ~n10885 & ~n10896;
  assign n10898 = ~n10884 & ~n10897;
  assign n10899 = ~n10883 & ~n10898;
  assign n10900 = ~n10882 & ~n10899;
  assign n10901 = ~n10881 & ~n10900;
  assign n10902 = ~n10880 & ~n10901;
  assign n10903 = ~pi200 & pi232;
  assign n10904 = pi199 & ~n10903;
  assign n10905 = ~n10902 & n10904;
  assign n10906 = pi231 & ~n10905;
  assign n10907 = ~n10902 & ~n10903;
  assign n10908 = ~pi199 & ~n10907;
  assign n10909 = ~n10906 & ~n10908;
  assign n10910 = pi200 & ~pi216;
  assign n10911 = ~pi201 & pi217;
  assign n10912 = pi201 & ~pi217;
  assign n10913 = ~pi202 & pi218;
  assign n10914 = pi202 & ~pi218;
  assign n10915 = ~pi203 & pi219;
  assign n10916 = pi203 & ~pi219;
  assign n10917 = ~pi205 & pi221;
  assign n10918 = pi206 & ~pi222;
  assign n10919 = ~n10917 & n10918;
  assign n10920 = pi205 & ~pi221;
  assign n10921 = pi204 & ~pi220;
  assign n10922 = ~n10920 & ~n10921;
  assign n10923 = ~n10919 & n10922;
  assign n10924 = ~pi204 & pi220;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926 = ~n10916 & ~n10925;
  assign n10927 = ~n10915 & ~n10926;
  assign n10928 = ~n10914 & ~n10927;
  assign n10929 = ~n10913 & ~n10928;
  assign n10930 = ~n10912 & ~n10929;
  assign n10931 = ~n10911 & ~n10930;
  assign n10932 = ~n10910 & ~n10931;
  assign n10933 = ~pi200 & pi216;
  assign n10934 = pi199 & ~n10933;
  assign n10935 = ~n10932 & n10934;
  assign n10936 = pi215 & ~n10935;
  assign n10937 = ~n10932 & ~n10933;
  assign n10938 = ~pi199 & ~n10937;
  assign n10939 = ~n10936 & ~n10938;
  assign n10940 = pi200 & ~pi224;
  assign n10941 = ~pi201 & pi225;
  assign n10942 = pi201 & ~pi225;
  assign n10943 = ~pi202 & pi226;
  assign n10944 = pi202 & ~pi226;
  assign n10945 = ~pi203 & pi227;
  assign n10946 = pi203 & ~pi227;
  assign n10947 = ~pi205 & pi229;
  assign n10948 = pi206 & ~pi230;
  assign n10949 = ~n10947 & n10948;
  assign n10950 = pi205 & ~pi229;
  assign n10951 = pi204 & ~pi228;
  assign n10952 = ~n10950 & ~n10951;
  assign n10953 = ~n10949 & n10952;
  assign n10954 = ~pi204 & pi228;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = ~n10946 & ~n10955;
  assign n10957 = ~n10945 & ~n10956;
  assign n10958 = ~n10944 & ~n10957;
  assign n10959 = ~n10943 & ~n10958;
  assign n10960 = ~n10942 & ~n10959;
  assign n10961 = ~n10941 & ~n10960;
  assign n10962 = ~n10940 & ~n10961;
  assign n10963 = ~pi200 & pi224;
  assign n10964 = pi199 & ~n10963;
  assign n10965 = ~n10962 & n10964;
  assign n10966 = pi223 & ~n10965;
  assign n10967 = ~n10962 & ~n10963;
  assign n10968 = ~pi199 & ~n10967;
  assign n10969 = ~n10966 & ~n10968;
  assign n10970 = ~n10939 & ~n10969;
  assign n10971 = ~n10909 & n10970;
  assign n10972 = ~n6371 & ~n7277;
  assign n10973 = n6181 & n10972;
  assign n10974 = ~n4578 & ~n5436;
  assign n10975 = n5732 & n10974;
  assign n10976 = n10973 & n10975;
  assign n10977 = ~n7385 & ~n8732;
  assign n10978 = ~n8820 & n10977;
  assign n10979 = ~n10818 & n10978;
  assign n10980 = n10976 & n10979;
  assign n10981 = ~n7358 & ~n8705;
  assign n10982 = ~n8793 & n10981;
  assign n10983 = ~n6344 & ~n7240;
  assign n10984 = n6740 & n10983;
  assign n10985 = ~n4551 & ~n5409;
  assign n10986 = n5757 & n10985;
  assign n10987 = n10984 & n10986;
  assign n10988 = n10982 & n10987;
  assign n10989 = ~n598 & ~n969;
  assign n10990 = ~n1145 & ~n2177;
  assign n10991 = n10989 & n10990;
  assign n10992 = n5718 & n10991;
  assign n10993 = ~n3256 & ~n3316;
  assign n10994 = ~n2455 & ~n2694;
  assign n10995 = n10993 & n10994;
  assign n10996 = n9873 & n10995;
  assign n10997 = n10992 & n10996;
  assign n10998 = n3861 & n10997;
  assign n10999 = n10988 & n10998;
  assign n11000 = ~n1172 & n10999;
  assign n11001 = ~n996 & n11000;
  assign n11002 = ~n2306 & n11001;
  assign n11003 = ~n500 & n11002;
  assign n11004 = ~n532 & ~n626;
  assign n11005 = n11003 & n11004;
  assign n11006 = ~n3283 & ~n3343;
  assign n11007 = ~n2482 & ~n2721;
  assign n11008 = n11006 & n11007;
  assign n11009 = n7601 & n11008;
  assign n11010 = n11005 & n11009;
  assign n11011 = n10980 & n11010;
  assign n11012 = n10971 & n11011;
  assign n11013 = pi200 & ~pi264;
  assign n11014 = ~pi201 & pi265;
  assign n11015 = pi201 & ~pi265;
  assign n11016 = ~pi202 & pi266;
  assign n11017 = pi202 & ~pi266;
  assign n11018 = ~pi203 & pi267;
  assign n11019 = pi203 & ~pi267;
  assign n11020 = ~pi204 & pi268;
  assign n11021 = pi204 & ~pi268;
  assign n11022 = pi206 & ~pi270;
  assign n11023 = pi205 & ~pi269;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = ~pi205 & pi269;
  assign n11026 = ~n11024 & ~n11025;
  assign n11027 = ~n11021 & ~n11026;
  assign n11028 = ~n11020 & ~n11027;
  assign n11029 = ~n11019 & ~n11028;
  assign n11030 = ~n11018 & ~n11029;
  assign n11031 = ~n11017 & ~n11030;
  assign n11032 = ~n11016 & ~n11031;
  assign n11033 = ~n11015 & ~n11032;
  assign n11034 = ~n11014 & ~n11033;
  assign n11035 = ~n11013 & ~n11034;
  assign n11036 = ~pi200 & pi264;
  assign n11037 = pi199 & ~n11036;
  assign n11038 = ~n11035 & n11037;
  assign n11039 = pi263 & ~n11038;
  assign n11040 = ~n11035 & ~n11036;
  assign n11041 = ~pi199 & ~n11040;
  assign n11042 = ~n11039 & ~n11041;
  assign n11043 = pi200 & ~pi256;
  assign n11044 = ~pi201 & pi257;
  assign n11045 = pi201 & ~pi257;
  assign n11046 = ~pi202 & pi258;
  assign n11047 = pi202 & ~pi258;
  assign n11048 = ~pi203 & pi259;
  assign n11049 = pi203 & ~pi259;
  assign n11050 = ~pi204 & pi260;
  assign n11051 = pi204 & ~pi260;
  assign n11052 = pi206 & ~pi262;
  assign n11053 = pi205 & ~pi261;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = ~pi205 & pi261;
  assign n11056 = ~n11054 & ~n11055;
  assign n11057 = ~n11051 & ~n11056;
  assign n11058 = ~n11050 & ~n11057;
  assign n11059 = ~n11049 & ~n11058;
  assign n11060 = ~n11048 & ~n11059;
  assign n11061 = ~n11047 & ~n11060;
  assign n11062 = ~n11046 & ~n11061;
  assign n11063 = ~n11045 & ~n11062;
  assign n11064 = ~n11044 & ~n11063;
  assign n11065 = ~n11043 & ~n11064;
  assign n11066 = ~pi200 & pi256;
  assign n11067 = pi199 & ~n11066;
  assign n11068 = ~n11065 & n11067;
  assign n11069 = pi255 & ~n11068;
  assign n11070 = ~n11065 & ~n11066;
  assign n11071 = ~pi199 & ~n11070;
  assign n11072 = ~n11069 & ~n11071;
  assign n11073 = ~n11042 & ~n11072;
  assign n11074 = pi200 & ~pi248;
  assign n11075 = ~pi201 & pi249;
  assign n11076 = pi201 & ~pi249;
  assign n11077 = ~pi202 & pi250;
  assign n11078 = pi202 & ~pi250;
  assign n11079 = ~pi203 & pi251;
  assign n11080 = pi203 & ~pi251;
  assign n11081 = ~pi204 & pi252;
  assign n11082 = pi204 & ~pi252;
  assign n11083 = pi206 & ~pi254;
  assign n11084 = pi205 & ~pi253;
  assign n11085 = ~n11083 & ~n11084;
  assign n11086 = ~pi205 & pi253;
  assign n11087 = ~n11085 & ~n11086;
  assign n11088 = ~n11082 & ~n11087;
  assign n11089 = ~n11081 & ~n11088;
  assign n11090 = ~n11080 & ~n11089;
  assign n11091 = ~n11079 & ~n11090;
  assign n11092 = ~n11078 & ~n11091;
  assign n11093 = ~n11077 & ~n11092;
  assign n11094 = ~n11076 & ~n11093;
  assign n11095 = ~n11075 & ~n11094;
  assign n11096 = ~n11074 & ~n11095;
  assign n11097 = ~pi200 & pi248;
  assign n11098 = pi199 & ~n11097;
  assign n11099 = ~n11096 & n11098;
  assign n11100 = pi247 & ~n11099;
  assign n11101 = ~n11096 & ~n11097;
  assign n11102 = ~pi199 & ~n11101;
  assign n11103 = ~n11100 & ~n11102;
  assign n11104 = pi200 & ~pi240;
  assign n11105 = ~pi201 & pi241;
  assign n11106 = pi201 & ~pi241;
  assign n11107 = ~pi202 & pi242;
  assign n11108 = pi202 & ~pi242;
  assign n11109 = ~pi203 & pi243;
  assign n11110 = pi203 & ~pi243;
  assign n11111 = ~pi204 & pi244;
  assign n11112 = pi204 & ~pi244;
  assign n11113 = pi206 & ~pi246;
  assign n11114 = pi205 & ~pi245;
  assign n11115 = ~n11113 & ~n11114;
  assign n11116 = ~pi205 & pi245;
  assign n11117 = ~n11115 & ~n11116;
  assign n11118 = ~n11112 & ~n11117;
  assign n11119 = ~n11111 & ~n11118;
  assign n11120 = ~n11110 & ~n11119;
  assign n11121 = ~n11109 & ~n11120;
  assign n11122 = ~n11108 & ~n11121;
  assign n11123 = ~n11107 & ~n11122;
  assign n11124 = ~n11106 & ~n11123;
  assign n11125 = ~n11105 & ~n11124;
  assign n11126 = ~n11104 & ~n11125;
  assign n11127 = ~pi200 & pi240;
  assign n11128 = pi199 & ~n11127;
  assign n11129 = ~n11126 & n11128;
  assign n11130 = pi239 & ~n11129;
  assign n11131 = ~n11126 & ~n11127;
  assign n11132 = ~pi199 & ~n11131;
  assign n11133 = ~n11130 & ~n11132;
  assign n11134 = ~n11103 & ~n11133;
  assign n11135 = n11073 & n11134;
  assign n11136 = ~n2080 & ~n2205;
  assign n11137 = n3822 & n11136;
  assign n11138 = n4787 & n11137;
  assign n11139 = pi200 & ~pi272;
  assign n11140 = ~pi201 & pi273;
  assign n11141 = pi201 & ~pi273;
  assign n11142 = ~pi202 & pi274;
  assign n11143 = pi202 & ~pi274;
  assign n11144 = ~pi203 & pi275;
  assign n11145 = pi203 & ~pi275;
  assign n11146 = ~pi204 & pi276;
  assign n11147 = pi204 & ~pi276;
  assign n11148 = pi206 & ~pi278;
  assign n11149 = pi205 & ~pi277;
  assign n11150 = ~n11148 & ~n11149;
  assign n11151 = ~pi205 & pi277;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n11147 & ~n11152;
  assign n11154 = ~n11146 & ~n11153;
  assign n11155 = ~n11145 & ~n11154;
  assign n11156 = ~n11144 & ~n11155;
  assign n11157 = ~n11143 & ~n11156;
  assign n11158 = ~n11142 & ~n11157;
  assign n11159 = ~n11141 & ~n11158;
  assign n11160 = ~n11140 & ~n11159;
  assign n11161 = ~n11139 & ~n11160;
  assign n11162 = ~pi200 & pi272;
  assign n11163 = pi199 & ~n11162;
  assign n11164 = ~n11161 & n11163;
  assign n11165 = pi271 & ~n11164;
  assign n11166 = ~n11161 & ~n11162;
  assign n11167 = ~pi199 & ~n11166;
  assign n11168 = ~n11165 & ~n11167;
  assign n11169 = n9592 & n9654;
  assign n11170 = ~n11168 & n11169;
  assign n11171 = n11138 & n11170;
  assign n11172 = n11135 & n11171;
  assign n11173 = n11012 & n11172;
  assign n11174 = ~n7236 & n11173;
  assign n11175 = ~n6137 & n11174;
  assign n11176 = n6193 & n11175;
  assign n11177 = n6134 & n11176;
  assign n11178 = ~n8867 & n11177;
  assign n11179 = ~n7235 & n11178;
  assign n11180 = n7296 & n11179;
  assign n11181 = n7231 & n11180;
  assign n11182 = ~n10027 & n11181;
  assign n11183 = ~n8866 & n11182;
  assign n11184 = n8898 & n11183;
  assign n11185 = n8863 & n11184;
  assign n11186 = ~n10026 & n11185;
  assign n11187 = n10072 & n11186;
  assign n11188 = n10021 & n11187;
  assign n11189 = ~n10879 & ~n11188;
  assign n11190 = ~n10787 & n11189;
  assign n11191 = n9654 & ~n10074;
  assign n11192 = ~n2453 & ~n3066;
  assign n11193 = ~n3983 & n11192;
  assign n11194 = ~n4024 & n11193;
  assign n11195 = ~n4999 & n11194;
  assign n11196 = ~n5827 & n11195;
  assign n11197 = ~n6893 & n11196;
  assign n11198 = ~n7890 & n11197;
  assign n11199 = ~n9131 & n11198;
  assign n11200 = ~n11191 & ~n11199;
  assign n11201 = ~n3524 & ~n3940;
  assign n11202 = ~n4001 & n11201;
  assign n11203 = ~n5043 & n11202;
  assign n11204 = ~n5943 & n11203;
  assign n11205 = ~n6951 & n11204;
  assign n11206 = ~n8037 & n11205;
  assign n11207 = ~n9200 & n11206;
  assign n11208 = ~n1649 & ~n2242;
  assign n11209 = ~n3095 & n11208;
  assign n11210 = ~n3997 & n11209;
  assign n11211 = ~n4837 & n11210;
  assign n11212 = ~n5822 & n11211;
  assign n11213 = ~n6820 & n11212;
  assign n11214 = ~n7785 & n11213;
  assign n11215 = ~n9027 & n11214;
  assign n11216 = ~n10245 & n11215;
  assign n11217 = ~n11207 & ~n11216;
  assign n11218 = n11200 & n11217;
  assign n11219 = n9718 & ~n9913;
  assign n11220 = n9624 & n11219;
  assign n11221 = n9856 & n11220;
  assign n11222 = ~n9929 & n11221;
  assign n11223 = ~n10416 & n11222;
  assign n11224 = ~n10622 & n11223;
  assign n11225 = n10564 & n11224;
  assign n11226 = ~n10713 & ~n10780;
  assign n11227 = n11225 & n11226;
  assign n11228 = n11218 & n11227;
  assign n11229 = ~n6461 & ~n6784;
  assign n11230 = ~n7158 & n11229;
  assign n11231 = ~n8250 & n11230;
  assign n11232 = ~n9414 & n11231;
  assign n11233 = ~n1115 & ~n1372;
  assign n11234 = ~n2243 & n11233;
  assign n11235 = ~n3104 & n11234;
  assign n11236 = ~n3971 & n11235;
  assign n11237 = ~n4872 & n11236;
  assign n11238 = ~n5801 & n11237;
  assign n11239 = ~n6739 & n11238;
  assign n11240 = ~n7807 & n11239;
  assign n11241 = ~n8989 & n11240;
  assign n11242 = ~n10273 & n11241;
  assign n11243 = ~n8662 & ~n8834;
  assign n11244 = ~n10002 & n11243;
  assign n11245 = ~n11242 & ~n11244;
  assign n11246 = ~n11232 & n11245;
  assign n11247 = ~n4677 & ~n4817;
  assign n11248 = ~n4902 & n11247;
  assign n11249 = ~n6001 & n11248;
  assign n11250 = ~n7014 & n11249;
  assign n11251 = ~n8114 & n11250;
  assign n11252 = ~n9276 & n11251;
  assign n11253 = ~n5527 & ~n5808;
  assign n11254 = ~n6056 & n11253;
  assign n11255 = ~n7073 & n11254;
  assign n11256 = ~n8179 & n11255;
  assign n11257 = ~n9344 & n11256;
  assign n11258 = ~n11252 & ~n11257;
  assign n11259 = ~n7327 & ~n7869;
  assign n11260 = ~n8346 & n11259;
  assign n11261 = ~n9485 & n11260;
  assign n11262 = ~n8900 & ~n9533;
  assign n11263 = ~n11261 & ~n11262;
  assign n11264 = n11258 & n11263;
  assign n11265 = n11246 & n11264;
  assign n11266 = n11228 & n11265;
  assign n11267 = ~n9200 & n9954;
  assign n11268 = ~n10713 & ~n11267;
  assign n11269 = ~n9344 & n9998;
  assign n11270 = ~n9533 & n9931;
  assign n11271 = ~n11269 & ~n11270;
  assign n11272 = n11268 & n11271;
  assign n11273 = n8662 & ~n9929;
  assign n11274 = n9934 & n9938;
  assign n11275 = n9937 & n11274;
  assign n11276 = n8545 & n11275;
  assign n11277 = ~n8834 & n11276;
  assign n11278 = ~n11273 & n11277;
  assign n11279 = ~n10416 & n11278;
  assign n11280 = ~n10002 & n11279;
  assign n11281 = ~n10780 & n11280;
  assign n11282 = n10640 & n11281;
  assign n11283 = n11272 & n11282;
  assign n11284 = n9994 & ~n10245;
  assign n11285 = ~n9485 & n9973;
  assign n11286 = ~n9414 & n9985;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = ~n11284 & n11287;
  assign n11289 = n8426 & ~n10074;
  assign n11290 = ~n9276 & n9971;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = ~n9131 & n9982;
  assign n11293 = n9966 & ~n10273;
  assign n11294 = ~n11292 & ~n11293;
  assign n11295 = n11291 & n11294;
  assign n11296 = n11288 & n11295;
  assign n11297 = n11283 & n11296;
  assign n11298 = ~n11266 & ~n11297;
  assign n11299 = ~n9344 & n10075;
  assign n11300 = ~n9276 & n10076;
  assign n11301 = ~n11299 & ~n11300;
  assign n11302 = ~n9200 & n10078;
  assign n11303 = ~n9131 & n10079;
  assign n11304 = ~n11302 & ~n11303;
  assign n11305 = n11301 & n11304;
  assign n11306 = ~n9485 & n10086;
  assign n11307 = n10083 & ~n10245;
  assign n11308 = ~n11306 & ~n11307;
  assign n11309 = n10082 & ~n10273;
  assign n11310 = ~n9414 & n10085;
  assign n11311 = ~n11309 & ~n11310;
  assign n11312 = n11308 & n11311;
  assign n11313 = n9515 & ~n10416;
  assign n11314 = ~n10094 & n11313;
  assign n11315 = ~n10713 & n11314;
  assign n11316 = n10640 & n11315;
  assign n11317 = n11312 & n11316;
  assign n11318 = n11305 & n11317;
  assign n11319 = ~n10713 & ~n11262;
  assign n11320 = ~n10002 & n10027;
  assign n11321 = ~n9485 & n10012;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = n11319 & n11322;
  assign n11324 = ~n9654 & ~n9929;
  assign n11325 = ~n10416 & ~n11324;
  assign n11326 = ~n10074 & n11325;
  assign n11327 = ~n10780 & n11326;
  assign n11328 = n10640 & n11327;
  assign n11329 = n11323 & n11328;
  assign n11330 = ~n9200 & n10070;
  assign n11331 = n10060 & ~n10273;
  assign n11332 = n10010 & ~n10245;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = ~n11330 & n11333;
  assign n11335 = ~n9131 & n10019;
  assign n11336 = ~n9276 & n10026;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = ~n9414 & n10064;
  assign n11339 = ~n9344 & n10051;
  assign n11340 = ~n11338 & ~n11339;
  assign n11341 = n11337 & n11340;
  assign n11342 = n11334 & n11341;
  assign n11343 = n11329 & n11342;
  assign n11344 = ~n11318 & ~n11343;
  assign n11345 = n11298 & n11344;
  assign po173 = ~n11190 | ~n11345;
  assign n11347 = ~n10763 & ~po173;
  assign n11348 = pi018 & ~n8900;
  assign n11349 = ~n10416 & n11348;
  assign n11350 = ~n9533 & n11349;
  assign n11351 = ~n10764 & n11350;
  assign n11352 = n10770 & n11351;
  assign n11353 = n10640 & n11352;
  assign n11354 = n10786 & n11353;
  assign n11355 = ~n8397 & n10162;
  assign n11356 = ~n10416 & n11355;
  assign n11357 = ~n10094 & n11356;
  assign n11358 = ~n10713 & n11357;
  assign n11359 = n10640 & n11358;
  assign n11360 = n11312 & n11359;
  assign n11361 = n11305 & n11360;
  assign n11362 = ~n11354 & ~n11361;
  assign n11363 = ~n9592 & ~n9717;
  assign n11364 = ~n9562 & ~n9622;
  assign n11365 = n11363 & n11364;
  assign n11366 = pi019 & ~n9687;
  assign n11367 = ~n9913 & n11366;
  assign n11368 = n11365 & n11367;
  assign n11369 = n9856 & n11368;
  assign n11370 = ~n9929 & n11369;
  assign n11371 = ~n10416 & n11370;
  assign n11372 = ~n10622 & n11371;
  assign n11373 = n10564 & n11372;
  assign n11374 = n11226 & n11373;
  assign n11375 = n11218 & n11374;
  assign n11376 = n11265 & n11375;
  assign n11377 = ~n8455 & ~n8633;
  assign n11378 = n8604 & n11377;
  assign n11379 = n10170 & n11378;
  assign n11380 = n9942 & n11379;
  assign n11381 = ~n8834 & n11380;
  assign n11382 = ~n11273 & n11381;
  assign n11383 = ~n10416 & n11382;
  assign n11384 = ~n10002 & n11383;
  assign n11385 = ~n10780 & n11384;
  assign n11386 = n10640 & n11385;
  assign n11387 = n11272 & n11386;
  assign n11388 = n11296 & n11387;
  assign n11389 = ~n11376 & ~n11388;
  assign n11390 = n11362 & n11389;
  assign n11391 = ~n11343 & ~n11390;
  assign n11392 = pi020 & ~n11324;
  assign n11393 = ~n10416 & n11392;
  assign n11394 = ~n10074 & n11393;
  assign n11395 = ~n10780 & n11394;
  assign n11396 = n10640 & n11395;
  assign n11397 = n11323 & n11396;
  assign n11398 = n11342 & n11397;
  assign n11399 = ~n6314 & ~n7387;
  assign n11400 = ~n8705 & ~n8764;
  assign n11401 = n11399 & n11400;
  assign n11402 = n4796 & n10836;
  assign n11403 = n7242 & n11402;
  assign n11404 = n11401 & n11403;
  assign n11405 = pi022 & ~n501;
  assign n11406 = ~n504 & ~n628;
  assign n11407 = n5713 & n11406;
  assign n11408 = n11405 & n11407;
  assign n11409 = ~n2052 & ~n2114;
  assign n11410 = n2219 & n11409;
  assign n11411 = n4846 & n11410;
  assign n11412 = n10136 & n10846;
  assign n11413 = n11411 & n11412;
  assign n11414 = n11408 & n11413;
  assign n11415 = n11404 & n11414;
  assign n11416 = ~n1172 & n11415;
  assign n11417 = ~n996 & n11416;
  assign n11418 = ~n2306 & n11417;
  assign n11419 = ~n500 & n11418;
  assign n11420 = n10855 & n11419;
  assign n11421 = n10860 & n11420;
  assign n11422 = n10831 & n11421;
  assign n11423 = n10823 & n11422;
  assign n11424 = ~n7236 & n11423;
  assign n11425 = ~n6137 & n11424;
  assign n11426 = n6193 & n11425;
  assign n11427 = n6134 & n11426;
  assign n11428 = ~n8867 & n11427;
  assign n11429 = ~n7295 & n11428;
  assign n11430 = n7231 & n11429;
  assign n11431 = ~n10788 & n11430;
  assign n11432 = ~n6344 & ~n7358;
  assign n11433 = ~n8705 & ~n8793;
  assign n11434 = n11432 & n11433;
  assign n11435 = n4796 & n10985;
  assign n11436 = n7242 & n11435;
  assign n11437 = n11434 & n11436;
  assign n11438 = pi021 & ~n501;
  assign n11439 = ~n504 & ~n598;
  assign n11440 = n5713 & n11439;
  assign n11441 = n11438 & n11440;
  assign n11442 = ~n2052 & ~n2177;
  assign n11443 = n2219 & n11442;
  assign n11444 = n4846 & n11443;
  assign n11445 = n10136 & n10995;
  assign n11446 = n11444 & n11445;
  assign n11447 = n11441 & n11446;
  assign n11448 = n11437 & n11447;
  assign n11449 = ~n1172 & n11448;
  assign n11450 = ~n996 & n11449;
  assign n11451 = ~n2306 & n11450;
  assign n11452 = ~n500 & n11451;
  assign n11453 = n11004 & n11452;
  assign n11454 = n11009 & n11453;
  assign n11455 = n10980 & n11454;
  assign n11456 = n10971 & n11455;
  assign n11457 = n11172 & n11456;
  assign n11458 = ~n7236 & n11457;
  assign n11459 = ~n6137 & n11458;
  assign n11460 = n6193 & n11459;
  assign n11461 = n6134 & n11460;
  assign n11462 = ~n8867 & n11461;
  assign n11463 = ~n7295 & n11462;
  assign n11464 = n7231 & n11463;
  assign n11465 = ~n11431 & ~n11464;
  assign n11466 = ~n7235 & ~n7293;
  assign n11467 = ~n10027 & n11466;
  assign n11468 = ~n8866 & n11467;
  assign n11469 = n8898 & n11468;
  assign n11470 = n8863 & n11469;
  assign n11471 = ~n10026 & n11470;
  assign n11472 = ~n11465 & n11471;
  assign n11473 = n10072 & n11472;
  assign n11474 = n10021 & n11473;
  assign n11475 = ~n11398 & ~n11474;
  assign n11476 = ~n11391 & n11475;
  assign po011 = n11347 | ~n11476;
  assign n11478 = n10780 & ~n11318;
  assign n11479 = ~n11266 & n11324;
  assign n11480 = ~n11478 & ~n11479;
  assign n11481 = n843 & n1239;
  assign n11482 = n720 & n11481;
  assign n11483 = ~n1372 & n11482;
  assign n11484 = ~n2243 & n11483;
  assign n11485 = ~n3104 & n11484;
  assign n11486 = ~n3837 & n11485;
  assign n11487 = ~n3971 & n11486;
  assign n11488 = ~n4872 & n11487;
  assign n11489 = ~n5801 & n11488;
  assign n11490 = ~n6739 & n11489;
  assign n11491 = ~n7807 & n11490;
  assign n11492 = ~n8989 & n11491;
  assign n11493 = ~n10293 & n11492;
  assign n11494 = ~n10292 & n11493;
  assign n11495 = ~n10273 & n11494;
  assign n11496 = ~n10291 & n11495;
  assign n11497 = n10290 & n11496;
  assign n11498 = n10285 & n11497;
  assign n11499 = n10326 & n11498;
  assign n11500 = n11331 & ~n11499;
  assign n11501 = ~n10705 & n10713;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = n11480 & n11502;
  assign n11504 = n10547 & ~n10554;
  assign n11505 = n10622 & ~n10629;
  assign n11506 = n10452 & ~n10460;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 = ~n11504 & n11507;
  assign n11509 = ~n10787 & n11262;
  assign n11510 = ~n10400 & n10416;
  assign n11511 = ~n10074 & ~n11510;
  assign n11512 = ~n11343 & n11511;
  assign n11513 = ~n11509 & n11512;
  assign n11514 = n11508 & n11513;
  assign n11515 = n11503 & n11514;
  assign n11516 = ~n10741 & n11321;
  assign n11517 = ~n1679 & ~n2206;
  assign n11518 = n1741 & n11517;
  assign n11519 = n3088 & n11518;
  assign n11520 = n1619 & n11519;
  assign n11521 = ~n2242 & n11520;
  assign n11522 = ~n3095 & n11521;
  assign n11523 = ~n3997 & n11522;
  assign n11524 = ~n4003 & n11523;
  assign n11525 = ~n4837 & n11524;
  assign n11526 = ~n5822 & n11525;
  assign n11527 = ~n6820 & n11526;
  assign n11528 = ~n7785 & n11527;
  assign n11529 = ~n9027 & n11528;
  assign n11530 = ~n10342 & n11529;
  assign n11531 = ~n10341 & n11530;
  assign n11532 = ~n10245 & n11531;
  assign n11533 = ~n10340 & n11532;
  assign n11534 = n10339 & n11533;
  assign n11535 = n10334 & n11534;
  assign n11536 = n10372 & n11535;
  assign n11537 = n11332 & ~n11536;
  assign n11538 = ~n11516 & ~n11537;
  assign n11539 = ~n10667 & n11338;
  assign n11540 = ~n11297 & n11320;
  assign n11541 = ~n11539 & ~n11540;
  assign n11542 = n11538 & n11541;
  assign n11543 = ~n10523 & n11336;
  assign n11544 = ~n10278 & n11335;
  assign n11545 = ~n11543 & ~n11544;
  assign n11546 = ~n10445 & n11330;
  assign n11547 = ~n10594 & n11339;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = n11545 & n11548;
  assign n11550 = n11542 & n11549;
  assign n11551 = n11515 & n11550;
  assign n11552 = ~n11478 & ~n11501;
  assign n11553 = ~n10445 & n11207;
  assign n11554 = n11242 & ~n11499;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = n11552 & n11555;
  assign n11557 = n9592 & ~n11188;
  assign n11558 = n9562 & ~n10879;
  assign n11559 = ~n9793 & ~n9824;
  assign n11560 = ~n9854 & n11559;
  assign n11561 = ~n9622 & n9718;
  assign n11562 = ~n9763 & ~n9913;
  assign n11563 = n11561 & n11562;
  assign n11564 = n11560 & n11563;
  assign n11565 = ~n9929 & n11564;
  assign n11566 = ~n11558 & n11565;
  assign n11567 = ~n11557 & n11566;
  assign n11568 = ~n11510 & n11567;
  assign n11569 = ~n11266 & n11568;
  assign n11570 = ~n11509 & n11569;
  assign n11571 = n11508 & n11570;
  assign n11572 = n11556 & n11571;
  assign n11573 = n11216 & ~n11536;
  assign n11574 = n11191 & ~n11343;
  assign n11575 = ~n11573 & ~n11574;
  assign n11576 = ~n10741 & n11261;
  assign n11577 = ~n10278 & n11199;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = n11575 & n11578;
  assign n11580 = ~n10667 & n11232;
  assign n11581 = ~n10523 & n11252;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = n11244 & ~n11297;
  assign n11584 = ~n10594 & n11257;
  assign n11585 = ~n11583 & ~n11584;
  assign n11586 = n11582 & n11585;
  assign n11587 = n11579 & n11586;
  assign n11588 = n11572 & n11587;
  assign n11589 = n11262 & ~n11510;
  assign n11590 = ~n10787 & n11589;
  assign n11591 = ~n11478 & n11590;
  assign n11592 = ~n10445 & n10783;
  assign n11593 = ~n11501 & ~n11592;
  assign n11594 = n11591 & n11593;
  assign n11595 = n11508 & n11594;
  assign n11596 = ~n10594 & n10764;
  assign n11597 = n10782 & ~n11499;
  assign n11598 = ~n11596 & ~n11597;
  assign n11599 = n10775 & ~n11536;
  assign n11600 = n10779 & ~n11297;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = n11598 & n11601;
  assign n11603 = ~n10667 & n10768;
  assign n11604 = ~n10278 & n10776;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = ~n10741 & n10769;
  assign n11607 = ~n10523 & n10773;
  assign n11608 = ~n11606 & ~n11607;
  assign n11609 = n11605 & n11608;
  assign n11610 = n11602 & n11609;
  assign n11611 = n11595 & n11610;
  assign n11612 = n10206 & ~n11266;
  assign n11613 = n10225 & ~n11297;
  assign n11614 = ~n11612 & ~n11613;
  assign n11615 = n10193 & ~n10741;
  assign n11616 = n10251 & ~n10523;
  assign n11617 = ~n11615 & ~n11616;
  assign n11618 = n11614 & n11617;
  assign n11619 = n10200 & ~n10629;
  assign n11620 = n10201 & ~n10554;
  assign n11621 = n10199 & ~n10460;
  assign n11622 = ~n11620 & ~n11621;
  assign n11623 = ~n11619 & n11622;
  assign n11624 = n10274 & ~n11499;
  assign n11625 = n10205 & ~n10400;
  assign n11626 = n2512 & ~n10879;
  assign n11627 = n2483 & ~n11188;
  assign n11628 = ~n2424 & ~n2754;
  assign n11629 = n9136 & n11628;
  assign n11630 = n2633 & n11629;
  assign n11631 = ~n3066 & n11630;
  assign n11632 = ~n3983 & n11631;
  assign n11633 = ~n4003 & n11632;
  assign n11634 = ~n4024 & n11633;
  assign n11635 = ~n4999 & n11634;
  assign n11636 = ~n5827 & n11635;
  assign n11637 = ~n6893 & n11636;
  assign n11638 = ~n7890 & n11637;
  assign n11639 = ~n9131 & n11638;
  assign n11640 = ~n11627 & n11639;
  assign n11641 = ~n11626 & n11640;
  assign n11642 = ~n11625 & n11641;
  assign n11643 = ~n10278 & n11642;
  assign n11644 = ~n11624 & n11643;
  assign n11645 = n11623 & n11644;
  assign n11646 = n11618 & n11645;
  assign n11647 = n10246 & ~n11536;
  assign n11648 = n10195 & ~n11343;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = n10253 & ~n11318;
  assign n11651 = n10250 & ~n10787;
  assign n11652 = ~n11650 & ~n11651;
  assign n11653 = n11649 & n11652;
  assign n11654 = n10204 & ~n10594;
  assign n11655 = n10196 & ~n10445;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = n10192 & ~n10667;
  assign n11658 = n10247 & ~n10705;
  assign n11659 = ~n11657 & ~n11658;
  assign n11660 = n11656 & n11659;
  assign n11661 = n11653 & n11660;
  assign n11662 = n11646 & n11661;
  assign n11663 = n10314 & ~n11297;
  assign n11664 = n10315 & ~n10741;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = n10319 & ~n10667;
  assign n11667 = n10282 & ~n10445;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = n11665 & n11668;
  assign n11670 = n10287 & ~n10629;
  assign n11671 = n10288 & ~n10554;
  assign n11672 = n10286 & ~n10460;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = ~n11670 & n11673;
  assign n11675 = n10323 & ~n11536;
  assign n11676 = n10292 & ~n10400;
  assign n11677 = n627 & ~n11188;
  assign n11678 = n657 & ~n10879;
  assign n11679 = ~n688 & ~n841;
  assign n11680 = ~n718 & n11679;
  assign n11681 = n4920 & n4929;
  assign n11682 = n10294 & n11681;
  assign n11683 = n11680 & n11682;
  assign n11684 = ~n1372 & n11683;
  assign n11685 = ~n2243 & n11684;
  assign n11686 = ~n3104 & n11685;
  assign n11687 = ~n3971 & n11686;
  assign n11688 = ~n4003 & n11687;
  assign n11689 = ~n4872 & n11688;
  assign n11690 = ~n5801 & n11689;
  assign n11691 = ~n6739 & n11690;
  assign n11692 = ~n7807 & n11691;
  assign n11693 = ~n8989 & n11692;
  assign n11694 = ~n10273 & n11693;
  assign n11695 = ~n11678 & n11694;
  assign n11696 = ~n11677 & n11695;
  assign n11697 = ~n11676 & n11696;
  assign n11698 = ~n11499 & n11697;
  assign n11699 = ~n11675 & n11698;
  assign n11700 = n11674 & n11699;
  assign n11701 = n11669 & n11700;
  assign n11702 = n10293 & ~n11266;
  assign n11703 = n10291 & ~n11343;
  assign n11704 = ~n11702 & ~n11703;
  assign n11705 = n10322 & ~n11318;
  assign n11706 = n10283 & ~n10787;
  assign n11707 = ~n11705 & ~n11706;
  assign n11708 = n11704 & n11707;
  assign n11709 = n10320 & ~n10523;
  assign n11710 = ~n10278 & n10279;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = n10280 & ~n10594;
  assign n11713 = n10316 & ~n10705;
  assign n11714 = ~n11712 & ~n11713;
  assign n11715 = n11711 & n11714;
  assign n11716 = n11708 & n11715;
  assign n11717 = n11701 & n11716;
  assign n11718 = n10360 & ~n11297;
  assign n11719 = n10361 & ~n10741;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 = n10365 & ~n10667;
  assign n11722 = n10331 & ~n10445;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = n11720 & n11723;
  assign n11725 = n10336 & ~n10629;
  assign n11726 = n10337 & ~n10554;
  assign n11727 = n10335 & ~n10460;
  assign n11728 = ~n11726 & ~n11727;
  assign n11729 = ~n11725 & n11728;
  assign n11730 = n10369 & ~n11499;
  assign n11731 = n10341 & ~n10400;
  assign n11732 = n2206 & ~n11188;
  assign n11733 = n2143 & ~n10879;
  assign n11734 = pi003 & ~n2176;
  assign n11735 = n4955 & n11734;
  assign n11736 = n7909 & n11735;
  assign n11737 = ~n2242 & n11736;
  assign n11738 = ~n3095 & n11737;
  assign n11739 = ~n3997 & n11738;
  assign n11740 = ~n4003 & n11739;
  assign n11741 = ~n4837 & n11740;
  assign n11742 = ~n5822 & n11741;
  assign n11743 = ~n6820 & n11742;
  assign n11744 = ~n7785 & n11743;
  assign n11745 = ~n9027 & n11744;
  assign n11746 = ~n10245 & n11745;
  assign n11747 = ~n11733 & n11746;
  assign n11748 = ~n11732 & n11747;
  assign n11749 = ~n11731 & n11748;
  assign n11750 = ~n11536 & n11749;
  assign n11751 = ~n11730 & n11750;
  assign n11752 = n11729 & n11751;
  assign n11753 = n11724 & n11752;
  assign n11754 = n10342 & ~n11266;
  assign n11755 = n10340 & ~n11343;
  assign n11756 = ~n11754 & ~n11755;
  assign n11757 = n10368 & ~n11318;
  assign n11758 = n10332 & ~n10787;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = n11756 & n11759;
  assign n11761 = n10366 & ~n10523;
  assign n11762 = ~n10278 & n10328;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 = n10329 & ~n10594;
  assign n11765 = n10362 & ~n10705;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = n11763 & n11766;
  assign n11768 = n11760 & n11767;
  assign n11769 = n11753 & n11768;
  assign n11770 = ~n11717 & ~n11769;
  assign n11771 = ~n11662 & n11770;
  assign n11772 = n7973 & n9115;
  assign n11773 = ~n3066 & n11772;
  assign n11774 = ~n3983 & n11773;
  assign n11775 = ~n4003 & n11774;
  assign n11776 = ~n4024 & n11775;
  assign n11777 = ~n4999 & n11776;
  assign n11778 = ~n5827 & n11777;
  assign n11779 = ~n6893 & n11778;
  assign n11780 = ~n7890 & n11779;
  assign n11781 = ~n9131 & n11780;
  assign n11782 = ~n11627 & n11781;
  assign n11783 = ~n11626 & n11782;
  assign n11784 = ~n11625 & n11783;
  assign n11785 = ~n10278 & n11784;
  assign n11786 = ~n11624 & n11785;
  assign n11787 = n11623 & n11786;
  assign n11788 = n11618 & n11787;
  assign n11789 = n11661 & n11788;
  assign n11790 = n10398 & ~n11499;
  assign n11791 = n10395 & ~n10400;
  assign n11792 = ~n11790 & n11791;
  assign n11793 = ~n10278 & n10394;
  assign n11794 = n10397 & ~n11536;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = n11792 & n11795;
  assign n11797 = ~n11789 & ~n11796;
  assign n11798 = ~n11771 & n11797;
  assign n11799 = n10417 & ~n11266;
  assign n11800 = n10432 & ~n11297;
  assign n11801 = ~n11799 & ~n11800;
  assign n11802 = n10437 & ~n10741;
  assign n11803 = n10438 & ~n10523;
  assign n11804 = ~n11802 & ~n11803;
  assign n11805 = n11801 & n11804;
  assign n11806 = n10410 & ~n10460;
  assign n11807 = n10411 & ~n10629;
  assign n11808 = n10412 & ~n10554;
  assign n11809 = ~n11807 & ~n11808;
  assign n11810 = ~n11806 & n11809;
  assign n11811 = n10433 & ~n11536;
  assign n11812 = n3373 & ~n10879;
  assign n11813 = n3344 & ~n11188;
  assign n11814 = ~n3403 & ~n3650;
  assign n11815 = n3621 & n11814;
  assign n11816 = n3800 & n11815;
  assign n11817 = ~n3940 & n11816;
  assign n11818 = ~n4001 & n11817;
  assign n11819 = ~n5043 & n11818;
  assign n11820 = ~n5943 & n11819;
  assign n11821 = ~n6951 & n11820;
  assign n11822 = ~n8037 & n11821;
  assign n11823 = ~n9200 & n11822;
  assign n11824 = ~n11813 & n11823;
  assign n11825 = ~n11812 & n11824;
  assign n11826 = ~n11510 & n11825;
  assign n11827 = ~n10445 & n11826;
  assign n11828 = ~n11811 & n11827;
  assign n11829 = n11810 & n11828;
  assign n11830 = n11805 & n11829;
  assign n11831 = n10403 & ~n10787;
  assign n11832 = n10440 & ~n11499;
  assign n11833 = ~n11831 & ~n11832;
  assign n11834 = n10441 & ~n11318;
  assign n11835 = n10434 & ~n10705;
  assign n11836 = ~n11834 & ~n11835;
  assign n11837 = n11833 & n11836;
  assign n11838 = n10404 & ~n10594;
  assign n11839 = ~n10278 & n10407;
  assign n11840 = ~n11838 & ~n11839;
  assign n11841 = n10415 & ~n10667;
  assign n11842 = n10406 & ~n11343;
  assign n11843 = ~n11841 & ~n11842;
  assign n11844 = n11840 & n11843;
  assign n11845 = n11837 & n11844;
  assign n11846 = n11830 & n11845;
  assign n11847 = ~n10400 & n10446;
  assign n11848 = ~n11790 & n11847;
  assign n11849 = n11795 & n11848;
  assign n11850 = ~n11846 & ~n11849;
  assign n11851 = ~n11798 & n11850;
  assign n11852 = ~n10278 & n10456;
  assign n11853 = n11506 & ~n11510;
  assign n11854 = ~n11852 & n11853;
  assign n11855 = ~n10445 & n10455;
  assign n11856 = n10457 & ~n11536;
  assign n11857 = n10451 & ~n11499;
  assign n11858 = ~n11856 & ~n11857;
  assign n11859 = ~n11855 & n11858;
  assign n11860 = n11854 & n11859;
  assign n11861 = ~n3403 & n4103;
  assign n11862 = n5062 & n10461;
  assign n11863 = n11861 & n11862;
  assign n11864 = ~n3940 & n11863;
  assign n11865 = ~n4001 & n11864;
  assign n11866 = ~n5043 & n11865;
  assign n11867 = ~n5943 & n11866;
  assign n11868 = ~n6951 & n11867;
  assign n11869 = ~n8037 & n11868;
  assign n11870 = ~n9200 & n11869;
  assign n11871 = ~n11813 & n11870;
  assign n11872 = ~n11812 & n11871;
  assign n11873 = ~n11510 & n11872;
  assign n11874 = ~n10445 & n11873;
  assign n11875 = ~n11811 & n11874;
  assign n11876 = n11810 & n11875;
  assign n11877 = n11805 & n11876;
  assign n11878 = n11845 & n11877;
  assign n11879 = ~n11860 & ~n11878;
  assign n11880 = ~n11851 & n11879;
  assign n11881 = ~n10460 & n10480;
  assign n11882 = ~n11510 & n11881;
  assign n11883 = ~n11852 & n11882;
  assign n11884 = n11859 & n11883;
  assign n11885 = n10510 & ~n11297;
  assign n11886 = n10516 & ~n10594;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = n10496 & ~n11266;
  assign n11889 = n10515 & ~n10741;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = n11887 & n11890;
  assign n11892 = n10491 & ~n10554;
  assign n11893 = n10492 & ~n10629;
  assign n11894 = ~n11506 & ~n11893;
  assign n11895 = ~n11892 & n11894;
  assign n11896 = n10519 & ~n11499;
  assign n11897 = n4579 & ~n11188;
  assign n11898 = n4608 & ~n10879;
  assign n11899 = n7030 & n8119;
  assign n11900 = ~n4817 & n11899;
  assign n11901 = ~n4902 & n11900;
  assign n11902 = ~n6001 & n11901;
  assign n11903 = ~n7014 & n11902;
  assign n11904 = ~n8114 & n11903;
  assign n11905 = ~n9276 & n11904;
  assign n11906 = ~n11898 & n11905;
  assign n11907 = ~n11897 & n11906;
  assign n11908 = ~n11510 & n11907;
  assign n11909 = ~n10523 & n11908;
  assign n11910 = ~n11896 & n11909;
  assign n11911 = n11895 & n11910;
  assign n11912 = n11891 & n11911;
  assign n11913 = n10511 & ~n11536;
  assign n11914 = n10487 & ~n11343;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 = n10512 & ~n11318;
  assign n11917 = n10484 & ~n10787;
  assign n11918 = ~n11916 & ~n11917;
  assign n11919 = n11915 & n11918;
  assign n11920 = ~n10445 & n10495;
  assign n11921 = ~n10278 & n10488;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = n10485 & ~n10667;
  assign n11924 = n10518 & ~n10705;
  assign n11925 = ~n11923 & ~n11924;
  assign n11926 = n11922 & n11925;
  assign n11927 = n11919 & n11926;
  assign n11928 = n11912 & n11927;
  assign n11929 = ~n11884 & ~n11928;
  assign n11930 = ~n11880 & n11929;
  assign n11931 = ~n4341 & n8095;
  assign n11932 = n5085 & n10526;
  assign n11933 = n11931 & n11932;
  assign n11934 = ~n4817 & n11933;
  assign n11935 = ~n4902 & n11934;
  assign n11936 = ~n6001 & n11935;
  assign n11937 = ~n7014 & n11936;
  assign n11938 = ~n8114 & n11937;
  assign n11939 = ~n9276 & n11938;
  assign n11940 = ~n11898 & n11939;
  assign n11941 = ~n11897 & n11940;
  assign n11942 = ~n11510 & n11941;
  assign n11943 = ~n10523 & n11942;
  assign n11944 = ~n11896 & n11943;
  assign n11945 = n11895 & n11944;
  assign n11946 = n11891 & n11945;
  assign n11947 = n11927 & n11946;
  assign n11948 = n10544 & ~n11536;
  assign n11949 = ~n10523 & n10551;
  assign n11950 = n10542 & ~n11499;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = ~n11948 & n11951;
  assign n11953 = n11504 & ~n11510;
  assign n11954 = ~n11506 & n11953;
  assign n11955 = ~n10445 & n10550;
  assign n11956 = ~n10278 & n10543;
  assign n11957 = ~n11955 & ~n11956;
  assign n11958 = n11954 & n11957;
  assign n11959 = n11952 & n11958;
  assign n11960 = ~n11947 & ~n11959;
  assign n11961 = ~n11930 & n11960;
  assign n11962 = n10581 & ~n11297;
  assign n11963 = n10586 & ~n10741;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = n10582 & ~n11536;
  assign n11966 = ~n10445 & n10567;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = n11964 & n11967;
  assign n11969 = n10565 & ~n10629;
  assign n11970 = ~n11504 & ~n11506;
  assign n11971 = ~n11969 & n11970;
  assign n11972 = n10590 & ~n11499;
  assign n11973 = n5437 & ~n11188;
  assign n11974 = n5289 & ~n10879;
  assign n11975 = ~n5230 & ~n5408;
  assign n11976 = n5379 & n11975;
  assign n11977 = n5688 & n11976;
  assign n11978 = ~n5808 & n11977;
  assign n11979 = ~n6056 & n11978;
  assign n11980 = ~n7073 & n11979;
  assign n11981 = ~n8179 & n11980;
  assign n11982 = ~n9344 & n11981;
  assign n11983 = ~n11974 & n11982;
  assign n11984 = ~n11973 & n11983;
  assign n11985 = ~n11510 & n11984;
  assign n11986 = ~n10594 & n11985;
  assign n11987 = ~n11972 & n11986;
  assign n11988 = n11971 & n11987;
  assign n11989 = n11968 & n11988;
  assign n11990 = n10560 & ~n11343;
  assign n11991 = n10568 & ~n11266;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = n10557 & ~n10787;
  assign n11994 = n10583 & ~n11318;
  assign n11995 = ~n11993 & ~n11994;
  assign n11996 = n11992 & n11995;
  assign n11997 = ~n10523 & n10587;
  assign n11998 = ~n10278 & n10561;
  assign n11999 = ~n11997 & ~n11998;
  assign n12000 = n10558 & ~n10667;
  assign n12001 = n10589 & ~n10705;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = n11999 & n12002;
  assign n12004 = n11996 & n12003;
  assign n12005 = n11989 & n12004;
  assign n12006 = ~n10554 & n10595;
  assign n12007 = ~n11510 & n12006;
  assign n12008 = ~n11506 & n12007;
  assign n12009 = n11957 & n12008;
  assign n12010 = n11952 & n12009;
  assign n12011 = ~n12005 & ~n12010;
  assign n12012 = ~n11961 & n12011;
  assign n12013 = ~n5230 & n6065;
  assign n12014 = n8190 & n12013;
  assign n12015 = ~n5808 & n12014;
  assign n12016 = ~n6056 & n12015;
  assign n12017 = ~n7073 & n12016;
  assign n12018 = ~n8179 & n12017;
  assign n12019 = ~n9344 & n12018;
  assign n12020 = ~n11974 & n12019;
  assign n12021 = ~n11973 & n12020;
  assign n12022 = ~n11510 & n12021;
  assign n12023 = ~n10594 & n12022;
  assign n12024 = ~n11972 & n12023;
  assign n12025 = n11971 & n12024;
  assign n12026 = n11968 & n12025;
  assign n12027 = n12004 & n12026;
  assign n12028 = ~n10278 & n10615;
  assign n12029 = ~n10594 & n10625;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = n10619 & ~n11536;
  assign n12032 = n10618 & ~n11499;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = n12030 & n12033;
  assign n12035 = n11505 & ~n11510;
  assign n12036 = n11970 & n12035;
  assign n12037 = ~n10523 & n10616;
  assign n12038 = ~n10445 & n10626;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = n12036 & n12039;
  assign n12041 = n12034 & n12040;
  assign n12042 = ~n12027 & ~n12041;
  assign n12043 = ~n12012 & n12042;
  assign n12044 = n10654 & ~n11297;
  assign n12045 = n10659 & ~n10741;
  assign n12046 = ~n12044 & ~n12045;
  assign n12047 = n10642 & ~n11266;
  assign n12048 = ~n10445 & n10660;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = n12046 & n12049;
  assign n12051 = n10655 & ~n11536;
  assign n12052 = n6372 & ~n11188;
  assign n12053 = n6342 & ~n10879;
  assign n12054 = ~n6313 & ~n6401;
  assign n12055 = n6614 & n12054;
  assign n12056 = n8236 & n12055;
  assign n12057 = ~n6784 & n12056;
  assign n12058 = ~n7158 & n12057;
  assign n12059 = ~n8250 & n12058;
  assign n12060 = ~n9414 & n12059;
  assign n12061 = ~n12053 & n12060;
  assign n12062 = ~n12052 & n12061;
  assign n12063 = ~n11510 & n12062;
  assign n12064 = ~n10667 & n12063;
  assign n12065 = ~n12051 & n12064;
  assign n12066 = n11508 & n12065;
  assign n12067 = n12050 & n12066;
  assign n12068 = n10635 & ~n11343;
  assign n12069 = n10663 & ~n11499;
  assign n12070 = ~n12068 & ~n12069;
  assign n12071 = n10656 & ~n11318;
  assign n12072 = n10633 & ~n10787;
  assign n12073 = ~n12071 & ~n12072;
  assign n12074 = n12070 & n12073;
  assign n12075 = ~n10523 & n10641;
  assign n12076 = ~n10278 & n10636;
  assign n12077 = ~n12075 & ~n12076;
  assign n12078 = ~n10594 & n10632;
  assign n12079 = n10662 & ~n10705;
  assign n12080 = ~n12078 & ~n12079;
  assign n12081 = n12077 & n12080;
  assign n12082 = n12074 & n12081;
  assign n12083 = n12067 & n12082;
  assign n12084 = ~n10629 & n10668;
  assign n12085 = ~n11510 & n12084;
  assign n12086 = n11970 & n12085;
  assign n12087 = n12039 & n12086;
  assign n12088 = n12034 & n12087;
  assign n12089 = ~n12083 & ~n12088;
  assign n12090 = ~n12043 & n12089;
  assign n12091 = n7177 & n10675;
  assign n12092 = n8261 & n12091;
  assign n12093 = ~n6784 & n12092;
  assign n12094 = ~n7158 & n12093;
  assign n12095 = ~n8250 & n12094;
  assign n12096 = ~n9414 & n12095;
  assign n12097 = ~n12053 & n12096;
  assign n12098 = ~n12052 & n12097;
  assign n12099 = ~n11510 & n12098;
  assign n12100 = ~n10667 & n12099;
  assign n12101 = ~n12051 & n12100;
  assign n12102 = n11508 & n12101;
  assign n12103 = n12050 & n12102;
  assign n12104 = n12082 & n12103;
  assign n12105 = ~n10523 & n10693;
  assign n12106 = n10700 & ~n11536;
  assign n12107 = ~n12105 & ~n12106;
  assign n12108 = n10696 & ~n11499;
  assign n12109 = ~n10445 & n10701;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = n12107 & n12110;
  assign n12112 = ~n10667 & n10689;
  assign n12113 = n10713 & ~n11510;
  assign n12114 = ~n10705 & n12113;
  assign n12115 = ~n12112 & n12114;
  assign n12116 = ~n10594 & n10690;
  assign n12117 = ~n10278 & n10692;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = n12115 & n12118;
  assign n12120 = n11508 & n12119;
  assign n12121 = n12111 & n12120;
  assign n12122 = n10737 & ~n11536;
  assign n12123 = n10728 & ~n11297;
  assign n12124 = ~n12122 & ~n12123;
  assign n12125 = ~n10667 & n10729;
  assign n12126 = n10714 & ~n11266;
  assign n12127 = ~n12125 & ~n12126;
  assign n12128 = n12124 & n12127;
  assign n12129 = n7386 & ~n11188;
  assign n12130 = n7415 & ~n10879;
  assign n12131 = n7476 & n10715;
  assign n12132 = n7753 & n12131;
  assign n12133 = ~n7869 & n12132;
  assign n12134 = ~n8346 & n12133;
  assign n12135 = ~n9485 & n12134;
  assign n12136 = ~n12130 & n12135;
  assign n12137 = ~n12129 & n12136;
  assign n12138 = ~n11510 & n12137;
  assign n12139 = ~n10741 & n12138;
  assign n12140 = ~n11501 & n12139;
  assign n12141 = n11508 & n12140;
  assign n12142 = n12128 & n12141;
  assign n12143 = n10733 & ~n10787;
  assign n12144 = n10710 & ~n11343;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = n10730 & ~n11499;
  assign n12147 = n10736 & ~n11318;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = n12145 & n12148;
  assign n12150 = ~n10445 & n10706;
  assign n12151 = ~n10523 & n10707;
  assign n12152 = ~n12150 & ~n12151;
  assign n12153 = ~n10278 & n10734;
  assign n12154 = ~n10594 & n10709;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = n12152 & n12155;
  assign n12157 = n12149 & n12156;
  assign n12158 = n12142 & n12157;
  assign n12159 = ~n12121 & ~n12158;
  assign n12160 = ~n12104 & n12159;
  assign n12161 = ~n12090 & n12160;
  assign n12162 = ~n10667 & n11310;
  assign n12163 = ~n10445 & n11302;
  assign n12164 = ~n12162 & ~n12163;
  assign n12165 = ~n10278 & n11303;
  assign n12166 = ~n10523 & n11300;
  assign n12167 = ~n12165 & ~n12166;
  assign n12168 = n12164 & n12167;
  assign n12169 = ~n10741 & n11306;
  assign n12170 = ~n10594 & n11299;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = n11309 & ~n11499;
  assign n12173 = n11307 & ~n11536;
  assign n12174 = ~n12172 & ~n12173;
  assign n12175 = n12171 & n12174;
  assign n12176 = n10780 & ~n11510;
  assign n12177 = ~n11318 & n12176;
  assign n12178 = ~n11501 & n12177;
  assign n12179 = n11508 & n12178;
  assign n12180 = n12175 & n12179;
  assign n12181 = n12168 & n12180;
  assign n12182 = ~n7356 & n8364;
  assign n12183 = n8361 & n12182;
  assign n12184 = ~n7869 & n12183;
  assign n12185 = ~n8346 & n12184;
  assign n12186 = ~n9485 & n12185;
  assign n12187 = ~n12130 & n12186;
  assign n12188 = ~n12129 & n12187;
  assign n12189 = ~n11510 & n12188;
  assign n12190 = ~n10741 & n12189;
  assign n12191 = ~n11501 & n12190;
  assign n12192 = n11508 & n12191;
  assign n12193 = n12128 & n12192;
  assign n12194 = n12157 & n12193;
  assign n12195 = ~n9453 & n10745;
  assign n12196 = ~n11510 & n12195;
  assign n12197 = ~n10705 & n12196;
  assign n12198 = ~n12112 & n12197;
  assign n12199 = n12118 & n12198;
  assign n12200 = n11508 & n12199;
  assign n12201 = n12111 & n12200;
  assign n12202 = ~n12194 & ~n12201;
  assign n12203 = ~n12181 & n12202;
  assign n12204 = ~n12161 & n12203;
  assign n12205 = ~n10278 & n11292;
  assign n12206 = ~n11501 & ~n12205;
  assign n12207 = ~n10741 & n11285;
  assign n12208 = ~n11266 & n11273;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = n12206 & n12209;
  assign n12211 = n8821 & ~n11188;
  assign n12212 = n8792 & ~n10879;
  assign n12213 = ~n8574 & ~n8762;
  assign n12214 = n9934 & n12213;
  assign n12215 = n8545 & n12214;
  assign n12216 = ~n8834 & n12215;
  assign n12217 = ~n10002 & n12216;
  assign n12218 = ~n12212 & n12217;
  assign n12219 = ~n12211 & n12218;
  assign n12220 = ~n11510 & n12219;
  assign n12221 = ~n11297 & n12220;
  assign n12222 = ~n11478 & n12221;
  assign n12223 = n11508 & n12222;
  assign n12224 = n12210 & n12223;
  assign n12225 = n11289 & ~n11343;
  assign n12226 = n11293 & ~n11499;
  assign n12227 = ~n12225 & ~n12226;
  assign n12228 = n11284 & ~n11536;
  assign n12229 = ~n10787 & n11270;
  assign n12230 = ~n12228 & ~n12229;
  assign n12231 = n12227 & n12230;
  assign n12232 = ~n10594 & n11269;
  assign n12233 = ~n10667 & n11286;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = ~n10445 & n11267;
  assign n12236 = ~n10523 & n11290;
  assign n12237 = ~n12235 & ~n12236;
  assign n12238 = n12234 & n12237;
  assign n12239 = n12231 & n12238;
  assign n12240 = n12224 & n12239;
  assign n12241 = ~pi016 & ~po161;
  assign n12242 = ~n8397 & n12241;
  assign n12243 = ~n10094 & n12242;
  assign n12244 = ~n11510 & n12243;
  assign n12245 = ~n11318 & n12244;
  assign n12246 = ~n11501 & n12245;
  assign n12247 = n11508 & n12246;
  assign n12248 = n12175 & n12247;
  assign n12249 = n12168 & n12248;
  assign n12250 = ~n12240 & ~n12249;
  assign n12251 = ~n12204 & n12250;
  assign n12252 = n10169 & n11378;
  assign n12253 = n9942 & n12252;
  assign n12254 = ~n8834 & n12253;
  assign n12255 = ~n10002 & n12254;
  assign n12256 = ~n12212 & n12255;
  assign n12257 = ~n12211 & n12256;
  assign n12258 = ~n11510 & n12257;
  assign n12259 = ~n11297 & n12258;
  assign n12260 = ~n11478 & n12259;
  assign n12261 = n11508 & n12260;
  assign n12262 = n12210 & n12261;
  assign n12263 = n12239 & n12262;
  assign n12264 = ~n12251 & ~n12263;
  assign n12265 = ~n11611 & ~n12264;
  assign n12266 = ~n9533 & n11348;
  assign n12267 = ~n11510 & n12266;
  assign n12268 = ~n10787 & n12267;
  assign n12269 = ~n11478 & n12268;
  assign n12270 = n11593 & n12269;
  assign n12271 = n11508 & n12270;
  assign n12272 = n11610 & n12271;
  assign n12273 = ~n12265 & ~n12272;
  assign n12274 = ~n11588 & ~n12273;
  assign n12275 = ~n9622 & ~n9717;
  assign n12276 = n11366 & n12275;
  assign n12277 = n11562 & n12276;
  assign n12278 = n11560 & n12277;
  assign n12279 = ~n9929 & n12278;
  assign n12280 = ~n11558 & n12279;
  assign n12281 = ~n11557 & n12280;
  assign n12282 = ~n11510 & n12281;
  assign n12283 = ~n11266 & n12282;
  assign n12284 = ~n11509 & n12283;
  assign n12285 = n11508 & n12284;
  assign n12286 = n11556 & n12285;
  assign n12287 = n11587 & n12286;
  assign n12288 = ~n12274 & ~n12287;
  assign n12289 = ~n11551 & ~n12288;
  assign n12290 = ~n627 & ~n1372;
  assign n12291 = ~n2243 & n12290;
  assign n12292 = ~n3104 & n12291;
  assign n12293 = ~n3971 & n12292;
  assign n12294 = ~n4872 & n12293;
  assign n12295 = ~n5801 & n12294;
  assign n12296 = ~n6739 & n12295;
  assign n12297 = ~n7807 & n12296;
  assign n12298 = ~n8989 & n12297;
  assign n12299 = ~n10273 & n12298;
  assign n12300 = ~n11499 & n12299;
  assign n12301 = ~n11501 & ~n12300;
  assign n12302 = ~n4579 & ~n4817;
  assign n12303 = ~n4902 & n12302;
  assign n12304 = ~n6001 & n12303;
  assign n12305 = ~n7014 & n12304;
  assign n12306 = ~n8114 & n12305;
  assign n12307 = ~n9276 & n12306;
  assign n12308 = ~n10523 & n12307;
  assign n12309 = ~n8821 & ~n8834;
  assign n12310 = ~n10002 & n12309;
  assign n12311 = ~n11297 & n12310;
  assign n12312 = ~n12308 & ~n12311;
  assign n12313 = n12301 & n12312;
  assign n12314 = n10818 & ~n10879;
  assign n12315 = ~n11072 & ~n11103;
  assign n12316 = ~n11133 & n12315;
  assign n12317 = ~n11042 & ~n11168;
  assign n12318 = n10971 & n12317;
  assign n12319 = n12316 & n12318;
  assign n12320 = ~n11188 & n12319;
  assign n12321 = ~n12314 & n12320;
  assign n12322 = ~n11510 & n12321;
  assign n12323 = ~n11505 & n12322;
  assign n12324 = n11970 & n12323;
  assign n12325 = ~n11478 & ~n11509;
  assign n12326 = n12324 & n12325;
  assign n12327 = n12313 & n12326;
  assign n12328 = ~n3344 & ~n3940;
  assign n12329 = ~n4001 & n12328;
  assign n12330 = ~n5043 & n12329;
  assign n12331 = ~n5943 & n12330;
  assign n12332 = ~n6951 & n12331;
  assign n12333 = ~n8037 & n12332;
  assign n12334 = ~n9200 & n12333;
  assign n12335 = ~n10445 & n12334;
  assign n12336 = ~n6372 & ~n6784;
  assign n12337 = ~n7158 & n12336;
  assign n12338 = ~n8250 & n12337;
  assign n12339 = ~n9414 & n12338;
  assign n12340 = ~n10667 & n12339;
  assign n12341 = ~n12335 & ~n12340;
  assign n12342 = ~n9592 & ~n9929;
  assign n12343 = ~n11266 & n12342;
  assign n12344 = ~n7386 & ~n7869;
  assign n12345 = ~n8346 & n12344;
  assign n12346 = ~n9485 & n12345;
  assign n12347 = ~n10741 & n12346;
  assign n12348 = ~n12343 & ~n12347;
  assign n12349 = n12341 & n12348;
  assign n12350 = ~n2483 & ~n3066;
  assign n12351 = ~n3983 & n12350;
  assign n12352 = ~n4024 & n12351;
  assign n12353 = ~n4999 & n12352;
  assign n12354 = ~n5827 & n12353;
  assign n12355 = ~n6893 & n12354;
  assign n12356 = ~n7890 & n12355;
  assign n12357 = ~n9131 & n12356;
  assign n12358 = ~n10278 & n12357;
  assign n12359 = ~n5437 & ~n5808;
  assign n12360 = ~n6056 & n12359;
  assign n12361 = ~n7073 & n12360;
  assign n12362 = ~n8179 & n12361;
  assign n12363 = ~n9344 & n12362;
  assign n12364 = ~n10594 & n12363;
  assign n12365 = ~n12358 & ~n12364;
  assign n12366 = ~n2206 & ~n2242;
  assign n12367 = ~n3095 & n12366;
  assign n12368 = ~n3997 & n12367;
  assign n12369 = ~n4837 & n12368;
  assign n12370 = ~n5822 & n12369;
  assign n12371 = ~n6820 & n12370;
  assign n12372 = ~n7785 & n12371;
  assign n12373 = ~n9027 & n12372;
  assign n12374 = ~n10245 & n12373;
  assign n12375 = ~n11536 & n12374;
  assign n12376 = ~n10074 & ~n11343;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = n12365 & n12377;
  assign n12379 = n12349 & n12378;
  assign n12380 = n12327 & n12379;
  assign n12381 = pi020 & ~n10074;
  assign n12382 = ~n11510 & n12381;
  assign n12383 = ~n11343 & n12382;
  assign n12384 = ~n11509 & n12383;
  assign n12385 = n11508 & n12384;
  assign n12386 = n11503 & n12385;
  assign n12387 = n11550 & n12386;
  assign n12388 = ~n12380 & ~n12387;
  assign n12389 = ~n12289 & n12388;
  assign n12390 = ~n11501 & ~n12376;
  assign n12391 = ~n657 & ~n1372;
  assign n12392 = ~n2243 & n12391;
  assign n12393 = ~n3104 & n12392;
  assign n12394 = ~n3971 & n12393;
  assign n12395 = ~n4872 & n12394;
  assign n12396 = ~n5801 & n12395;
  assign n12397 = ~n6739 & n12396;
  assign n12398 = ~n7807 & n12397;
  assign n12399 = ~n8989 & n12398;
  assign n12400 = ~n10273 & n12399;
  assign n12401 = ~n11499 & n12400;
  assign n12402 = ~n3373 & ~n3940;
  assign n12403 = ~n4001 & n12402;
  assign n12404 = ~n5043 & n12403;
  assign n12405 = ~n5943 & n12404;
  assign n12406 = ~n6951 & n12405;
  assign n12407 = ~n8037 & n12406;
  assign n12408 = ~n9200 & n12407;
  assign n12409 = ~n10445 & n12408;
  assign n12410 = ~n12401 & ~n12409;
  assign n12411 = n12390 & n12410;
  assign n12412 = ~n10818 & ~n11188;
  assign n12413 = ~n10879 & ~n12412;
  assign n12414 = ~n11510 & n12413;
  assign n12415 = ~n11505 & n12414;
  assign n12416 = n11970 & n12415;
  assign n12417 = n12325 & n12416;
  assign n12418 = n12411 & n12417;
  assign n12419 = ~n8792 & ~n8834;
  assign n12420 = ~n10002 & n12419;
  assign n12421 = ~n11297 & n12420;
  assign n12422 = ~n4608 & ~n4817;
  assign n12423 = ~n4902 & n12422;
  assign n12424 = ~n6001 & n12423;
  assign n12425 = ~n7014 & n12424;
  assign n12426 = ~n8114 & n12425;
  assign n12427 = ~n9276 & n12426;
  assign n12428 = ~n10523 & n12427;
  assign n12429 = ~n12421 & ~n12428;
  assign n12430 = ~n5289 & ~n5808;
  assign n12431 = ~n6056 & n12430;
  assign n12432 = ~n7073 & n12431;
  assign n12433 = ~n8179 & n12432;
  assign n12434 = ~n9344 & n12433;
  assign n12435 = ~n10594 & n12434;
  assign n12436 = ~n2512 & ~n3066;
  assign n12437 = ~n3983 & n12436;
  assign n12438 = ~n4024 & n12437;
  assign n12439 = ~n4999 & n12438;
  assign n12440 = ~n5827 & n12439;
  assign n12441 = ~n6893 & n12440;
  assign n12442 = ~n7890 & n12441;
  assign n12443 = ~n9131 & n12442;
  assign n12444 = ~n10278 & n12443;
  assign n12445 = ~n12435 & ~n12444;
  assign n12446 = n12429 & n12445;
  assign n12447 = ~n2143 & ~n2242;
  assign n12448 = ~n3095 & n12447;
  assign n12449 = ~n3997 & n12448;
  assign n12450 = ~n4837 & n12449;
  assign n12451 = ~n5822 & n12450;
  assign n12452 = ~n6820 & n12451;
  assign n12453 = ~n7785 & n12452;
  assign n12454 = ~n9027 & n12453;
  assign n12455 = ~n10245 & n12454;
  assign n12456 = ~n11536 & n12455;
  assign n12457 = ~n6342 & ~n6784;
  assign n12458 = ~n7158 & n12457;
  assign n12459 = ~n8250 & n12458;
  assign n12460 = ~n9414 & n12459;
  assign n12461 = ~n10667 & n12460;
  assign n12462 = ~n12456 & ~n12461;
  assign n12463 = ~n7415 & ~n7869;
  assign n12464 = ~n8346 & n12463;
  assign n12465 = ~n9485 & n12464;
  assign n12466 = ~n10741 & n12465;
  assign n12467 = n10788 & ~n11266;
  assign n12468 = ~n12466 & ~n12467;
  assign n12469 = n12462 & n12468;
  assign n12470 = n12446 & n12469;
  assign n12471 = n12418 & n12470;
  assign n12472 = ~pi021 & ~n10939;
  assign n12473 = ~n10909 & ~n10969;
  assign n12474 = n12472 & n12473;
  assign n12475 = n12317 & n12474;
  assign n12476 = n12316 & n12475;
  assign n12477 = ~n11188 & n12476;
  assign n12478 = ~n12314 & n12477;
  assign n12479 = ~n11510 & n12478;
  assign n12480 = ~n11505 & n12479;
  assign n12481 = n11970 & n12480;
  assign n12482 = n12325 & n12481;
  assign n12483 = n12313 & n12482;
  assign n12484 = n12379 & n12483;
  assign n12485 = ~n12471 & ~n12484;
  assign n12486 = ~n12389 & n12485;
  assign n12487 = pi022 & ~n10879;
  assign n12488 = ~n12412 & n12487;
  assign n12489 = ~n11510 & n12488;
  assign n12490 = ~n11505 & n12489;
  assign n12491 = n11970 & n12490;
  assign n12492 = n12325 & n12491;
  assign n12493 = n12411 & n12492;
  assign n12494 = n12470 & n12493;
  assign n12495 = ~n1463 & ~n9651;
  assign n12496 = ~n9619 & ~n9653;
  assign n12497 = n12495 & n12496;
  assign n12498 = ~n2110 & ~n2175;
  assign n12499 = n4786 & n12498;
  assign n12500 = n12497 & n12499;
  assign n12501 = ~pi216 & pi224;
  assign n12502 = pi216 & ~pi224;
  assign n12503 = ~pi217 & pi225;
  assign n12504 = pi217 & ~pi225;
  assign n12505 = ~pi218 & pi226;
  assign n12506 = pi218 & ~pi226;
  assign n12507 = ~pi219 & pi227;
  assign n12508 = pi219 & ~pi227;
  assign n12509 = ~pi221 & pi229;
  assign n12510 = pi222 & ~pi230;
  assign n12511 = ~n12509 & n12510;
  assign n12512 = pi221 & ~pi229;
  assign n12513 = pi220 & ~pi228;
  assign n12514 = ~n12512 & ~n12513;
  assign n12515 = ~n12511 & n12514;
  assign n12516 = ~pi220 & pi228;
  assign n12517 = ~n12515 & ~n12516;
  assign n12518 = ~n12508 & ~n12517;
  assign n12519 = ~n12507 & ~n12518;
  assign n12520 = ~n12506 & ~n12519;
  assign n12521 = ~n12505 & ~n12520;
  assign n12522 = ~n12504 & ~n12521;
  assign n12523 = ~n12503 & ~n12522;
  assign n12524 = ~n12502 & ~n12523;
  assign n12525 = ~n12501 & ~n12524;
  assign n12526 = ~pi215 & ~n12525;
  assign n12527 = pi215 & ~n12501;
  assign n12528 = ~n12524 & n12527;
  assign n12529 = pi223 & ~n12528;
  assign n12530 = ~n10968 & ~n12529;
  assign n12531 = ~n12526 & n12530;
  assign n12532 = ~n9621 & ~n10815;
  assign n12533 = ~n10817 & ~n10966;
  assign n12534 = n12532 & n12533;
  assign n12535 = n12531 & n12534;
  assign n12536 = n12500 & n12535;
  assign n12537 = ~n8761 & ~n8791;
  assign n12538 = n10824 & n12537;
  assign n12539 = ~n6492 & ~n7355;
  assign n12540 = n10826 & n12539;
  assign n12541 = n6182 & n12540;
  assign n12542 = n12538 & n12541;
  assign n12543 = ~n8734 & n11400;
  assign n12544 = ~n6314 & ~n6465;
  assign n12545 = ~n7328 & ~n7387;
  assign n12546 = n12544 & n12545;
  assign n12547 = n7242 & n12546;
  assign n12548 = n12543 & n12547;
  assign n12549 = ~n2635 & ~n3375;
  assign n12550 = ~n4283 & ~n5570;
  assign n12551 = n12549 & n12550;
  assign n12552 = n11402 & n12551;
  assign n12553 = n11412 & n12552;
  assign n12554 = ~n534 & ~n782;
  assign n12555 = n11406 & n12554;
  assign n12556 = pi024 & ~n501;
  assign n12557 = n5713 & n12556;
  assign n12558 = n12555 & n12557;
  assign n12559 = ~n1404 & ~n2082;
  assign n12560 = ~n1435 & ~n2114;
  assign n12561 = n12559 & n12560;
  assign n12562 = ~n2052 & ~n2147;
  assign n12563 = n2219 & n12562;
  assign n12564 = n12561 & n12563;
  assign n12565 = n12558 & n12564;
  assign n12566 = n12553 & n12565;
  assign n12567 = n12548 & n12566;
  assign n12568 = ~n1172 & n12567;
  assign n12569 = ~n996 & n12568;
  assign n12570 = ~n2306 & n12569;
  assign n12571 = ~n2662 & ~n2691;
  assign n12572 = n12570 & n12571;
  assign n12573 = n6677 & n12572;
  assign n12574 = ~n4310 & ~n4607;
  assign n12575 = ~n5288 & ~n5597;
  assign n12576 = n12574 & n12575;
  assign n12577 = ~n3372 & ~n3402;
  assign n12578 = ~n2511 & ~n3254;
  assign n12579 = n12577 & n12578;
  assign n12580 = n12576 & n12579;
  assign n12581 = n12573 & n12580;
  assign n12582 = ~n656 & ~n810;
  assign n12583 = n3821 & n12582;
  assign n12584 = n10821 & n12583;
  assign n12585 = n12581 & n12584;
  assign n12586 = n12542 & n12585;
  assign n12587 = n12536 & n12586;
  assign n12588 = ~n7236 & n12587;
  assign n12589 = ~n6137 & n12588;
  assign n12590 = n6193 & n12589;
  assign n12591 = n6134 & n12590;
  assign n12592 = ~n8867 & n12591;
  assign n12593 = ~n7295 & n12592;
  assign n12594 = n7231 & n12593;
  assign n12595 = ~n10788 & n12594;
  assign n12596 = ~n8575 & n11400;
  assign n12597 = ~n6314 & ~n6644;
  assign n12598 = ~n7387 & ~n7418;
  assign n12599 = n12597 & n12598;
  assign n12600 = n7242 & n12599;
  assign n12601 = n12596 & n12600;
  assign n12602 = ~n3345 & ~n3770;
  assign n12603 = n4795 & n12602;
  assign n12604 = n3810 & n10845;
  assign n12605 = n12603 & n12604;
  assign n12606 = ~n2726 & ~n3256;
  assign n12607 = ~n4313 & ~n5202;
  assign n12608 = n12606 & n12607;
  assign n12609 = n11402 & n12608;
  assign n12610 = n12605 & n12609;
  assign n12611 = ~n534 & ~n812;
  assign n12612 = n11406 & n12611;
  assign n12613 = pi023 & ~n501;
  assign n12614 = n5713 & n12613;
  assign n12615 = n12612 & n12614;
  assign n12616 = ~n1588 & ~n2082;
  assign n12617 = n12560 & n12616;
  assign n12618 = n2219 & n5717;
  assign n12619 = n12617 & n12618;
  assign n12620 = n12615 & n12619;
  assign n12621 = n12610 & n12620;
  assign n12622 = n12601 & n12621;
  assign n12623 = ~n1172 & n12622;
  assign n12624 = ~n996 & n12623;
  assign n12625 = ~n2306 & n12624;
  assign n12626 = ~n2691 & ~n2753;
  assign n12627 = n12625 & n12626;
  assign n12628 = ~n656 & ~n840;
  assign n12629 = n12627 & n12628;
  assign n12630 = n3823 & n12629;
  assign n12631 = ~n1616 & ~n9651;
  assign n12632 = n4786 & n12631;
  assign n12633 = n3808 & n10820;
  assign n12634 = n12632 & n12633;
  assign n12635 = n12630 & n12634;
  assign n12636 = ~n8602 & ~n8791;
  assign n12637 = n10824 & n12636;
  assign n12638 = ~n6671 & ~n7445;
  assign n12639 = n10826 & n12638;
  assign n12640 = n12637 & n12639;
  assign n12641 = ~n12526 & ~n12529;
  assign n12642 = pi216 & ~pi232;
  assign n12643 = ~pi217 & pi233;
  assign n12644 = pi217 & ~pi233;
  assign n12645 = ~pi218 & pi234;
  assign n12646 = pi218 & ~pi234;
  assign n12647 = ~pi219 & pi235;
  assign n12648 = pi219 & ~pi235;
  assign n12649 = ~pi221 & pi237;
  assign n12650 = pi222 & ~pi238;
  assign n12651 = ~n12649 & n12650;
  assign n12652 = pi221 & ~pi237;
  assign n12653 = pi220 & ~pi236;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~n12651 & n12654;
  assign n12656 = ~pi220 & pi236;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12648 & ~n12657;
  assign n12659 = ~n12647 & ~n12658;
  assign n12660 = ~n12646 & ~n12659;
  assign n12661 = ~n12645 & ~n12660;
  assign n12662 = ~n12644 & ~n12661;
  assign n12663 = ~n12643 & ~n12662;
  assign n12664 = ~n12642 & ~n12663;
  assign n12665 = ~pi216 & pi232;
  assign n12666 = pi215 & ~n12665;
  assign n12667 = ~n12664 & n12666;
  assign n12668 = pi231 & ~n12667;
  assign n12669 = ~n12664 & ~n12665;
  assign n12670 = ~pi215 & ~n12669;
  assign n12671 = ~n12668 & ~n12670;
  assign n12672 = ~n12641 & ~n12671;
  assign n12673 = n12640 & n12672;
  assign n12674 = ~n3372 & ~n3797;
  assign n12675 = n12578 & n12674;
  assign n12676 = n6677 & n12675;
  assign n12677 = ~n4340 & ~n4607;
  assign n12678 = ~n5229 & ~n5288;
  assign n12679 = n12677 & n12678;
  assign n12680 = n6182 & n12679;
  assign n12681 = n12676 & n12680;
  assign n12682 = n12673 & n12681;
  assign n12683 = n12635 & n12682;
  assign n12684 = pi216 & ~pi256;
  assign n12685 = ~pi217 & pi257;
  assign n12686 = pi217 & ~pi257;
  assign n12687 = ~pi218 & pi258;
  assign n12688 = pi218 & ~pi258;
  assign n12689 = ~pi219 & pi259;
  assign n12690 = pi219 & ~pi259;
  assign n12691 = ~pi220 & pi260;
  assign n12692 = pi220 & ~pi260;
  assign n12693 = pi222 & ~pi262;
  assign n12694 = pi221 & ~pi261;
  assign n12695 = ~n12693 & ~n12694;
  assign n12696 = ~pi221 & pi261;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = ~n12692 & ~n12697;
  assign n12699 = ~n12691 & ~n12698;
  assign n12700 = ~n12690 & ~n12699;
  assign n12701 = ~n12689 & ~n12700;
  assign n12702 = ~n12688 & ~n12701;
  assign n12703 = ~n12687 & ~n12702;
  assign n12704 = ~n12686 & ~n12703;
  assign n12705 = ~n12685 & ~n12704;
  assign n12706 = ~n12684 & ~n12705;
  assign n12707 = ~pi216 & pi256;
  assign n12708 = pi215 & ~n12707;
  assign n12709 = ~n12706 & n12708;
  assign n12710 = pi255 & ~n12709;
  assign n12711 = ~n12706 & ~n12707;
  assign n12712 = ~pi215 & ~n12711;
  assign n12713 = ~n12710 & ~n12712;
  assign n12714 = pi216 & ~pi272;
  assign n12715 = ~pi217 & pi273;
  assign n12716 = pi217 & ~pi273;
  assign n12717 = ~pi218 & pi274;
  assign n12718 = pi218 & ~pi274;
  assign n12719 = ~pi219 & pi275;
  assign n12720 = pi219 & ~pi275;
  assign n12721 = ~pi220 & pi276;
  assign n12722 = pi220 & ~pi276;
  assign n12723 = pi222 & ~pi278;
  assign n12724 = pi221 & ~pi277;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = ~pi221 & pi277;
  assign n12727 = ~n12725 & ~n12726;
  assign n12728 = ~n12722 & ~n12727;
  assign n12729 = ~n12721 & ~n12728;
  assign n12730 = ~n12720 & ~n12729;
  assign n12731 = ~n12719 & ~n12730;
  assign n12732 = ~n12718 & ~n12731;
  assign n12733 = ~n12717 & ~n12732;
  assign n12734 = ~n12716 & ~n12733;
  assign n12735 = ~n12715 & ~n12734;
  assign n12736 = ~n12714 & ~n12735;
  assign n12737 = ~pi216 & pi272;
  assign n12738 = pi215 & ~n12737;
  assign n12739 = ~n12736 & n12738;
  assign n12740 = pi271 & ~n12739;
  assign n12741 = ~n12736 & ~n12737;
  assign n12742 = ~pi215 & ~n12741;
  assign n12743 = ~n12740 & ~n12742;
  assign n12744 = pi216 & ~pi264;
  assign n12745 = ~pi217 & pi265;
  assign n12746 = pi217 & ~pi265;
  assign n12747 = ~pi218 & pi266;
  assign n12748 = pi218 & ~pi266;
  assign n12749 = ~pi219 & pi267;
  assign n12750 = pi219 & ~pi267;
  assign n12751 = ~pi220 & pi268;
  assign n12752 = pi220 & ~pi268;
  assign n12753 = pi222 & ~pi270;
  assign n12754 = pi221 & ~pi269;
  assign n12755 = ~n12753 & ~n12754;
  assign n12756 = ~pi221 & pi269;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = ~n12752 & ~n12757;
  assign n12759 = ~n12751 & ~n12758;
  assign n12760 = ~n12750 & ~n12759;
  assign n12761 = ~n12749 & ~n12760;
  assign n12762 = ~n12748 & ~n12761;
  assign n12763 = ~n12747 & ~n12762;
  assign n12764 = ~n12746 & ~n12763;
  assign n12765 = ~n12745 & ~n12764;
  assign n12766 = ~n12744 & ~n12765;
  assign n12767 = ~pi216 & pi264;
  assign n12768 = pi215 & ~n12767;
  assign n12769 = ~n12766 & n12768;
  assign n12770 = pi263 & ~n12769;
  assign n12771 = ~n12766 & ~n12767;
  assign n12772 = ~pi215 & ~n12771;
  assign n12773 = ~n12770 & ~n12772;
  assign n12774 = ~n12743 & ~n12773;
  assign n12775 = ~n12713 & n12774;
  assign n12776 = ~n10817 & ~n10936;
  assign n12777 = ~n10938 & n12776;
  assign n12778 = ~n9653 & ~n9684;
  assign n12779 = ~n9686 & ~n10815;
  assign n12780 = n12778 & n12779;
  assign n12781 = n12777 & n12780;
  assign n12782 = pi216 & ~pi240;
  assign n12783 = ~pi217 & pi241;
  assign n12784 = pi217 & ~pi241;
  assign n12785 = ~pi218 & pi242;
  assign n12786 = pi218 & ~pi242;
  assign n12787 = ~pi219 & pi243;
  assign n12788 = pi219 & ~pi243;
  assign n12789 = ~pi220 & pi244;
  assign n12790 = pi220 & ~pi244;
  assign n12791 = pi222 & ~pi246;
  assign n12792 = pi221 & ~pi245;
  assign n12793 = ~n12791 & ~n12792;
  assign n12794 = ~pi221 & pi245;
  assign n12795 = ~n12793 & ~n12794;
  assign n12796 = ~n12790 & ~n12795;
  assign n12797 = ~n12789 & ~n12796;
  assign n12798 = ~n12788 & ~n12797;
  assign n12799 = ~n12787 & ~n12798;
  assign n12800 = ~n12786 & ~n12799;
  assign n12801 = ~n12785 & ~n12800;
  assign n12802 = ~n12784 & ~n12801;
  assign n12803 = ~n12783 & ~n12802;
  assign n12804 = ~n12782 & ~n12803;
  assign n12805 = ~pi216 & pi240;
  assign n12806 = pi215 & ~n12805;
  assign n12807 = ~n12804 & n12806;
  assign n12808 = pi239 & ~n12807;
  assign n12809 = ~n12804 & ~n12805;
  assign n12810 = ~pi215 & ~n12809;
  assign n12811 = ~n12808 & ~n12810;
  assign n12812 = pi216 & ~pi248;
  assign n12813 = ~pi217 & pi249;
  assign n12814 = pi217 & ~pi249;
  assign n12815 = ~pi218 & pi250;
  assign n12816 = pi218 & ~pi250;
  assign n12817 = ~pi219 & pi251;
  assign n12818 = pi219 & ~pi251;
  assign n12819 = ~pi220 & pi252;
  assign n12820 = pi220 & ~pi252;
  assign n12821 = pi222 & ~pi254;
  assign n12822 = pi221 & ~pi253;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = ~pi221 & pi253;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = ~n12820 & ~n12825;
  assign n12827 = ~n12819 & ~n12826;
  assign n12828 = ~n12818 & ~n12827;
  assign n12829 = ~n12817 & ~n12828;
  assign n12830 = ~n12816 & ~n12829;
  assign n12831 = ~n12815 & ~n12830;
  assign n12832 = ~n12814 & ~n12831;
  assign n12833 = ~n12813 & ~n12832;
  assign n12834 = ~n12812 & ~n12833;
  assign n12835 = ~pi216 & pi248;
  assign n12836 = pi215 & ~n12835;
  assign n12837 = ~n12834 & n12836;
  assign n12838 = pi247 & ~n12837;
  assign n12839 = ~n12834 & ~n12835;
  assign n12840 = ~pi215 & ~n12839;
  assign n12841 = ~n12838 & ~n12840;
  assign n12842 = ~n12811 & ~n12841;
  assign n12843 = n12781 & n12842;
  assign n12844 = n12775 & n12843;
  assign n12845 = n12683 & n12844;
  assign n12846 = ~n7236 & n12845;
  assign n12847 = ~n6137 & n12846;
  assign n12848 = n6193 & n12847;
  assign n12849 = n6134 & n12848;
  assign n12850 = ~n8867 & n12849;
  assign n12851 = ~n7295 & n12850;
  assign n12852 = n7231 & n12851;
  assign n12853 = ~n10788 & n12852;
  assign n12854 = ~n12595 & ~n12853;
  assign n12855 = n11471 & ~n12854;
  assign n12856 = n10072 & n12855;
  assign n12857 = n10021 & n12856;
  assign n12858 = ~n12494 & ~n12857;
  assign po012 = n12486 | ~n12858;
  assign n12860 = n11504 & ~n11959;
  assign n12861 = n11510 & ~n11796;
  assign n12862 = ~n8575 & ~n8764;
  assign n12863 = n12598 & n12862;
  assign n12864 = n10836 & n12597;
  assign n12865 = n12608 & n12864;
  assign n12866 = n12863 & n12865;
  assign n12867 = n10845 & n12602;
  assign n12868 = n3942 & n12867;
  assign n12869 = n8870 & n12868;
  assign n12870 = n4847 & n12611;
  assign n12871 = n4798 & n12616;
  assign n12872 = ~n628 & ~n1145;
  assign n12873 = n11409 & n12872;
  assign n12874 = n12871 & n12873;
  assign n12875 = n12870 & n12874;
  assign n12876 = n12869 & n12875;
  assign n12877 = n12866 & n12876;
  assign n12878 = ~n1172 & n12877;
  assign n12879 = ~n996 & n12878;
  assign n12880 = ~n2306 & n12879;
  assign n12881 = n12626 & n12880;
  assign n12882 = n12628 & n12881;
  assign n12883 = n3823 & n12882;
  assign n12884 = n12634 & n12883;
  assign n12885 = n12682 & n12884;
  assign n12886 = n12844 & n12885;
  assign n12887 = ~n7236 & n12886;
  assign n12888 = ~n6137 & n12887;
  assign n12889 = n6193 & n12888;
  assign n12890 = n6134 & n12889;
  assign n12891 = ~n8867 & n12890;
  assign n12892 = ~n7235 & n12891;
  assign n12893 = n7296 & n12892;
  assign n12894 = n7231 & n12893;
  assign n12895 = ~n10027 & n12894;
  assign n12896 = ~n8866 & n12895;
  assign n12897 = n8898 & n12896;
  assign n12898 = n8863 & n12897;
  assign n12899 = ~n10788 & n12898;
  assign n12900 = ~n10026 & n12899;
  assign n12901 = n10072 & n12900;
  assign n12902 = n10021 & n12901;
  assign n12903 = ~n12641 & ~n12902;
  assign n12904 = ~n8734 & ~n8764;
  assign n12905 = n12545 & n12904;
  assign n12906 = n10836 & n12544;
  assign n12907 = n8869 & n12906;
  assign n12908 = n12905 & n12907;
  assign n12909 = n3859 & n5757;
  assign n12910 = n7812 & n12909;
  assign n12911 = ~n2484 & ~n3345;
  assign n12912 = n4849 & n12911;
  assign n12913 = n12551 & n12912;
  assign n12914 = n12910 & n12913;
  assign n12915 = n4847 & n12554;
  assign n12916 = ~n2082 & ~n2147;
  assign n12917 = n4798 & n12916;
  assign n12918 = n12873 & n12917;
  assign n12919 = n12915 & n12918;
  assign n12920 = n12914 & n12919;
  assign n12921 = n12908 & n12920;
  assign n12922 = ~n1172 & n12921;
  assign n12923 = ~n996 & n12922;
  assign n12924 = ~n2306 & n12923;
  assign n12925 = n12571 & n12924;
  assign n12926 = n6677 & n12925;
  assign n12927 = n12580 & n12926;
  assign n12928 = n12584 & n12927;
  assign n12929 = n12542 & n12928;
  assign n12930 = n12536 & n12929;
  assign n12931 = ~n7236 & n12930;
  assign n12932 = ~n6137 & n12931;
  assign n12933 = n6193 & n12932;
  assign n12934 = n6134 & n12933;
  assign n12935 = ~n8867 & n12934;
  assign n12936 = ~n7235 & n12935;
  assign n12937 = n7296 & n12936;
  assign n12938 = n7231 & n12937;
  assign n12939 = ~n10027 & n12938;
  assign n12940 = ~n8866 & n12939;
  assign n12941 = n8898 & n12940;
  assign n12942 = n8863 & n12941;
  assign n12943 = ~n10788 & n12942;
  assign n12944 = ~n10026 & n12943;
  assign n12945 = n10072 & n12944;
  assign n12946 = n10021 & n12945;
  assign n12947 = ~n12903 & ~n12946;
  assign n12948 = ~n12861 & n12947;
  assign n12949 = ~n12860 & n12948;
  assign n12950 = n11506 & ~n11860;
  assign n12951 = n11505 & ~n12041;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = n12949 & n12952;
  assign n12954 = ~n3403 & ~n3940;
  assign n12955 = ~n4001 & n12954;
  assign n12956 = ~n5043 & n12955;
  assign n12957 = ~n5943 & n12956;
  assign n12958 = ~n6951 & n12957;
  assign n12959 = ~n8037 & n12958;
  assign n12960 = ~n9200 & n12959;
  assign n12961 = ~n10445 & n12960;
  assign n12962 = ~n11846 & n12961;
  assign n12963 = ~n4311 & ~n4817;
  assign n12964 = ~n4902 & n12963;
  assign n12965 = ~n6001 & n12964;
  assign n12966 = ~n7014 & n12965;
  assign n12967 = ~n8114 & n12966;
  assign n12968 = ~n9276 & n12967;
  assign n12969 = ~n10523 & n12968;
  assign n12970 = ~n11928 & n12969;
  assign n12971 = ~n12962 & ~n12970;
  assign n12972 = ~n11551 & n12376;
  assign n12973 = n11478 & ~n12181;
  assign n12974 = ~n12972 & ~n12973;
  assign n12975 = n12971 & n12974;
  assign n12976 = n12953 & n12975;
  assign n12977 = ~n2663 & ~n3066;
  assign n12978 = ~n3983 & n12977;
  assign n12979 = ~n4024 & n12978;
  assign n12980 = ~n4999 & n12979;
  assign n12981 = ~n5827 & n12980;
  assign n12982 = ~n6893 & n12981;
  assign n12983 = ~n7890 & n12982;
  assign n12984 = ~n9131 & n12983;
  assign n12985 = ~n10278 & n12984;
  assign n12986 = ~n11662 & n12985;
  assign n12987 = ~n9622 & ~n9929;
  assign n12988 = ~n11266 & n12987;
  assign n12989 = ~n11588 & n12988;
  assign n12990 = ~n12986 & ~n12989;
  assign n12991 = ~n8762 & ~n8834;
  assign n12992 = ~n10002 & n12991;
  assign n12993 = ~n11297 & n12992;
  assign n12994 = ~n12240 & n12993;
  assign n12995 = ~n7356 & ~n7869;
  assign n12996 = ~n8346 & n12995;
  assign n12997 = ~n9485 & n12996;
  assign n12998 = ~n10741 & n12997;
  assign n12999 = ~n12158 & n12998;
  assign n13000 = ~n12994 & ~n12999;
  assign n13001 = n12990 & n13000;
  assign n13002 = ~n5598 & ~n5808;
  assign n13003 = ~n6056 & n13002;
  assign n13004 = ~n7073 & n13003;
  assign n13005 = ~n8179 & n13004;
  assign n13006 = ~n9344 & n13005;
  assign n13007 = ~n10594 & n13006;
  assign n13008 = ~n12005 & n13007;
  assign n13009 = ~n6493 & ~n6784;
  assign n13010 = ~n7158 & n13009;
  assign n13011 = ~n8250 & n13010;
  assign n13012 = ~n9414 & n13011;
  assign n13013 = ~n10667 & n13012;
  assign n13014 = ~n12083 & n13013;
  assign n13015 = ~n13008 & ~n13014;
  assign n13016 = ~n1679 & ~n2176;
  assign n13017 = n1741 & n13016;
  assign n13018 = n1619 & n13017;
  assign n13019 = ~n2242 & n13018;
  assign n13020 = ~n3095 & n13019;
  assign n13021 = ~n3997 & n13020;
  assign n13022 = ~n4003 & n13021;
  assign n13023 = ~n4837 & n13022;
  assign n13024 = ~n5822 & n13023;
  assign n13025 = ~n6820 & n13024;
  assign n13026 = ~n7785 & n13025;
  assign n13027 = ~n9027 & n13026;
  assign n13028 = ~n10245 & n13027;
  assign n13029 = ~n11733 & n13028;
  assign n13030 = ~n11732 & n13029;
  assign n13031 = ~n11731 & n13030;
  assign n13032 = ~n11536 & n13031;
  assign n13033 = ~n11730 & n13032;
  assign n13034 = n11729 & n13033;
  assign n13035 = n11724 & n13034;
  assign n13036 = n11768 & n13035;
  assign n13037 = ~n2176 & ~n2242;
  assign n13038 = ~n3095 & n13037;
  assign n13039 = ~n3997 & n13038;
  assign n13040 = ~n4837 & n13039;
  assign n13041 = ~n5822 & n13040;
  assign n13042 = ~n6820 & n13041;
  assign n13043 = ~n7785 & n13042;
  assign n13044 = ~n9027 & n13043;
  assign n13045 = ~n10245 & n13044;
  assign n13046 = ~n11536 & n13045;
  assign n13047 = ~n13036 & n13046;
  assign n13048 = ~n10969 & ~n11188;
  assign n13049 = ~n12380 & n13048;
  assign n13050 = ~n13047 & ~n13049;
  assign n13051 = n13015 & n13050;
  assign n13052 = n11501 & ~n12121;
  assign n13053 = n11509 & ~n11611;
  assign n13054 = ~n13052 & ~n13053;
  assign n13055 = ~n10879 & ~n12471;
  assign n13056 = n719 & n842;
  assign n13057 = n2272 & n13056;
  assign n13058 = ~n1372 & n13057;
  assign n13059 = ~n2243 & n13058;
  assign n13060 = ~n3104 & n13059;
  assign n13061 = ~n3837 & n13060;
  assign n13062 = ~n3971 & n13061;
  assign n13063 = ~n4872 & n13062;
  assign n13064 = ~n5801 & n13063;
  assign n13065 = ~n6739 & n13064;
  assign n13066 = ~n7807 & n13065;
  assign n13067 = ~n8989 & n13066;
  assign n13068 = ~n10273 & n13067;
  assign n13069 = ~n11678 & n13068;
  assign n13070 = ~n11677 & n13069;
  assign n13071 = ~n11676 & n13070;
  assign n13072 = ~n11499 & n13071;
  assign n13073 = ~n11675 & n13072;
  assign n13074 = n11674 & n13073;
  assign n13075 = n11669 & n13074;
  assign n13076 = n11716 & n13075;
  assign n13077 = ~n811 & ~n1372;
  assign n13078 = ~n2243 & n13077;
  assign n13079 = ~n3104 & n13078;
  assign n13080 = ~n3971 & n13079;
  assign n13081 = ~n4872 & n13080;
  assign n13082 = ~n5801 & n13081;
  assign n13083 = ~n6739 & n13082;
  assign n13084 = ~n7807 & n13083;
  assign n13085 = ~n8989 & n13084;
  assign n13086 = ~n10273 & n13085;
  assign n13087 = ~n11499 & n13086;
  assign n13088 = ~n13076 & n13087;
  assign n13089 = ~n13055 & ~n13088;
  assign n13090 = n13054 & n13089;
  assign n13091 = n13051 & n13090;
  assign n13092 = n13001 & n13091;
  assign n13093 = n12976 & n13092;
  assign n13094 = ~n12860 & ~n12950;
  assign n13095 = ~n12951 & n13094;
  assign n13096 = n8762 & ~n12946;
  assign n13097 = n8603 & ~n12902;
  assign n13098 = ~n8574 & ~n8633;
  assign n13099 = n8545 & n13098;
  assign n13100 = ~n8834 & n13099;
  assign n13101 = ~n10002 & n13100;
  assign n13102 = ~n13097 & n13101;
  assign n13103 = ~n13096 & n13102;
  assign n13104 = ~n11297 & n13103;
  assign n13105 = ~n12861 & n13104;
  assign n13106 = ~n12240 & n13105;
  assign n13107 = ~n12973 & n13106;
  assign n13108 = ~n11588 & n12208;
  assign n13109 = ~n13052 & ~n13108;
  assign n13110 = n13107 & n13109;
  assign n13111 = n13095 & n13110;
  assign n13112 = ~n12083 & n12233;
  assign n13113 = n12228 & ~n13036;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = n12212 & ~n12471;
  assign n13116 = n12211 & ~n12380;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = n13114 & n13117;
  assign n13119 = n12226 & ~n13076;
  assign n13120 = ~n11928 & n12236;
  assign n13121 = ~n13119 & ~n13120;
  assign n13122 = ~n11611 & n12229;
  assign n13123 = ~n11551 & n12225;
  assign n13124 = ~n13122 & ~n13123;
  assign n13125 = n13121 & n13124;
  assign n13126 = ~n11662 & n12205;
  assign n13127 = ~n12158 & n12207;
  assign n13128 = ~n13126 & ~n13127;
  assign n13129 = ~n11846 & n12235;
  assign n13130 = ~n12005 & n12232;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = n13128 & n13131;
  assign n13133 = n13125 & n13132;
  assign n13134 = n13118 & n13133;
  assign n13135 = n13111 & n13134;
  assign n13136 = n11621 & ~n11860;
  assign n13137 = n11619 & ~n12041;
  assign n13138 = n11620 & ~n11959;
  assign n13139 = ~n13137 & ~n13138;
  assign n13140 = ~n13136 & n13139;
  assign n13141 = n11627 & ~n12380;
  assign n13142 = n11625 & ~n11796;
  assign n13143 = n2663 & ~n12946;
  assign n13144 = n2754 & ~n12902;
  assign n13145 = ~n2424 & ~n2783;
  assign n13146 = n2632 & n13145;
  assign n13147 = n2573 & n13146;
  assign n13148 = ~n3066 & n13147;
  assign n13149 = ~n3983 & n13148;
  assign n13150 = ~n4003 & n13149;
  assign n13151 = ~n4024 & n13150;
  assign n13152 = ~n4999 & n13151;
  assign n13153 = ~n5827 & n13152;
  assign n13154 = ~n6893 & n13153;
  assign n13155 = ~n7890 & n13154;
  assign n13156 = ~n9131 & n13155;
  assign n13157 = ~n13144 & n13156;
  assign n13158 = ~n13143 & n13157;
  assign n13159 = ~n10278 & n13158;
  assign n13160 = ~n13142 & n13159;
  assign n13161 = ~n11662 & n13160;
  assign n13162 = ~n13141 & n13161;
  assign n13163 = n11657 & ~n12083;
  assign n13164 = n11624 & ~n13076;
  assign n13165 = ~n13163 & ~n13164;
  assign n13166 = n13162 & n13165;
  assign n13167 = n13140 & n13166;
  assign n13168 = n11615 & ~n12158;
  assign n13169 = n11650 & ~n12181;
  assign n13170 = ~n13168 & ~n13169;
  assign n13171 = ~n11551 & n11648;
  assign n13172 = n11658 & ~n12121;
  assign n13173 = ~n13171 & ~n13172;
  assign n13174 = n13170 & n13173;
  assign n13175 = n11613 & ~n12240;
  assign n13176 = n11626 & ~n12471;
  assign n13177 = ~n13175 & ~n13176;
  assign n13178 = n11655 & ~n11846;
  assign n13179 = ~n11588 & n11612;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = n13177 & n13180;
  assign n13182 = n11616 & ~n11928;
  assign n13183 = ~n11611 & n11651;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = n11654 & ~n12005;
  assign n13186 = n11647 & ~n13036;
  assign n13187 = ~n13185 & ~n13186;
  assign n13188 = n13184 & n13187;
  assign n13189 = n13181 & n13188;
  assign n13190 = n13174 & n13189;
  assign n13191 = n13167 & n13190;
  assign n13192 = n11672 & ~n11860;
  assign n13193 = n11670 & ~n12041;
  assign n13194 = n11671 & ~n11959;
  assign n13195 = ~n13193 & ~n13194;
  assign n13196 = ~n13192 & n13195;
  assign n13197 = ~n11611 & n11706;
  assign n13198 = n11676 & ~n11796;
  assign n13199 = n841 & ~n12902;
  assign n13200 = n811 & ~n12946;
  assign n13201 = ~n688 & ~n780;
  assign n13202 = ~n718 & n13201;
  assign n13203 = n10295 & n13202;
  assign n13204 = ~n1372 & n13203;
  assign n13205 = ~n2243 & n13204;
  assign n13206 = ~n3104 & n13205;
  assign n13207 = ~n3971 & n13206;
  assign n13208 = ~n4003 & n13207;
  assign n13209 = ~n4872 & n13208;
  assign n13210 = ~n5801 & n13209;
  assign n13211 = ~n6739 & n13210;
  assign n13212 = ~n7807 & n13211;
  assign n13213 = ~n8989 & n13212;
  assign n13214 = ~n10273 & n13213;
  assign n13215 = ~n13200 & n13214;
  assign n13216 = ~n13199 & n13215;
  assign n13217 = ~n11499 & n13216;
  assign n13218 = ~n13198 & n13217;
  assign n13219 = ~n13076 & n13218;
  assign n13220 = ~n13197 & n13219;
  assign n13221 = n11712 & ~n12005;
  assign n13222 = n11667 & ~n11846;
  assign n13223 = ~n13221 & ~n13222;
  assign n13224 = n13220 & n13223;
  assign n13225 = n13196 & n13224;
  assign n13226 = n11666 & ~n12083;
  assign n13227 = n11705 & ~n12181;
  assign n13228 = ~n13226 & ~n13227;
  assign n13229 = ~n11551 & n11703;
  assign n13230 = n11713 & ~n12121;
  assign n13231 = ~n13229 & ~n13230;
  assign n13232 = n13228 & n13231;
  assign n13233 = n11675 & ~n13036;
  assign n13234 = ~n11588 & n11702;
  assign n13235 = ~n13233 & ~n13234;
  assign n13236 = ~n11662 & n11710;
  assign n13237 = n11663 & ~n12240;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = n13235 & n13238;
  assign n13240 = n11678 & ~n12471;
  assign n13241 = n11677 & ~n12380;
  assign n13242 = ~n13240 & ~n13241;
  assign n13243 = n11709 & ~n11928;
  assign n13244 = n11664 & ~n12158;
  assign n13245 = ~n13243 & ~n13244;
  assign n13246 = n13242 & n13245;
  assign n13247 = n13239 & n13246;
  assign n13248 = n13232 & n13247;
  assign n13249 = n13225 & n13248;
  assign n13250 = n11727 & ~n11860;
  assign n13251 = n11725 & ~n12041;
  assign n13252 = n11726 & ~n11959;
  assign n13253 = ~n13251 & ~n13252;
  assign n13254 = ~n13250 & n13253;
  assign n13255 = n11733 & ~n12471;
  assign n13256 = n11731 & ~n11796;
  assign n13257 = n1617 & ~n12902;
  assign n13258 = n2176 & ~n12946;
  assign n13259 = n1557 & ~n1587;
  assign n13260 = pi003 & ~n1679;
  assign n13261 = n1741 & n13260;
  assign n13262 = n13259 & n13261;
  assign n13263 = ~n2242 & n13262;
  assign n13264 = ~n3095 & n13263;
  assign n13265 = ~n3997 & n13264;
  assign n13266 = ~n4003 & n13265;
  assign n13267 = ~n4837 & n13266;
  assign n13268 = ~n5822 & n13267;
  assign n13269 = ~n6820 & n13268;
  assign n13270 = ~n7785 & n13269;
  assign n13271 = ~n9027 & n13270;
  assign n13272 = ~n10245 & n13271;
  assign n13273 = ~n13258 & n13272;
  assign n13274 = ~n13257 & n13273;
  assign n13275 = ~n11536 & n13274;
  assign n13276 = ~n13256 & n13275;
  assign n13277 = ~n13036 & n13276;
  assign n13278 = ~n13255 & n13277;
  assign n13279 = n11732 & ~n12380;
  assign n13280 = n11764 & ~n12005;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = n13278 & n13281;
  assign n13283 = n13254 & n13282;
  assign n13284 = ~n11662 & n11762;
  assign n13285 = n11757 & ~n12181;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = ~n11551 & n11755;
  assign n13288 = n11765 & ~n12121;
  assign n13289 = ~n13287 & ~n13288;
  assign n13290 = n13286 & n13289;
  assign n13291 = n11761 & ~n11928;
  assign n13292 = n11722 & ~n11846;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = ~n11611 & n11758;
  assign n13295 = ~n11588 & n11754;
  assign n13296 = ~n13294 & ~n13295;
  assign n13297 = n13293 & n13296;
  assign n13298 = n11730 & ~n13076;
  assign n13299 = n11718 & ~n12240;
  assign n13300 = ~n13298 & ~n13299;
  assign n13301 = n11721 & ~n12083;
  assign n13302 = n11719 & ~n12158;
  assign n13303 = ~n13301 & ~n13302;
  assign n13304 = n13300 & n13303;
  assign n13305 = n13297 & n13304;
  assign n13306 = n13290 & n13305;
  assign n13307 = n13283 & n13306;
  assign n13308 = ~n13249 & ~n13307;
  assign n13309 = ~n13191 & n13308;
  assign n13310 = n11794 & ~n13036;
  assign n13311 = ~n11790 & ~n11793;
  assign n13312 = ~n11794 & n13311;
  assign n13313 = n11791 & ~n13312;
  assign n13314 = ~n13310 & n13313;
  assign n13315 = ~n11662 & n11793;
  assign n13316 = n11790 & ~n13076;
  assign n13317 = ~n13315 & ~n13316;
  assign n13318 = n13314 & n13317;
  assign n13319 = ~n2783 & n3852;
  assign n13320 = n9134 & n13319;
  assign n13321 = ~n3066 & n13320;
  assign n13322 = ~n3983 & n13321;
  assign n13323 = ~n4003 & n13322;
  assign n13324 = ~n4024 & n13323;
  assign n13325 = ~n4999 & n13324;
  assign n13326 = ~n5827 & n13325;
  assign n13327 = ~n6893 & n13326;
  assign n13328 = ~n7890 & n13327;
  assign n13329 = ~n9131 & n13328;
  assign n13330 = ~n13144 & n13329;
  assign n13331 = ~n13143 & n13330;
  assign n13332 = ~n10278 & n13331;
  assign n13333 = ~n13142 & n13332;
  assign n13334 = ~n11662 & n13333;
  assign n13335 = ~n13141 & n13334;
  assign n13336 = n13165 & n13335;
  assign n13337 = n13140 & n13336;
  assign n13338 = n13190 & n13337;
  assign n13339 = ~n13318 & ~n13338;
  assign n13340 = ~n13309 & n13339;
  assign n13341 = n11808 & ~n11959;
  assign n13342 = n11806 & ~n11860;
  assign n13343 = n11807 & ~n12041;
  assign n13344 = ~n13342 & ~n13343;
  assign n13345 = ~n13341 & n13344;
  assign n13346 = n11841 & ~n12083;
  assign n13347 = n3798 & ~n12902;
  assign n13348 = n3403 & ~n12946;
  assign n13349 = ~n3591 & ~n3769;
  assign n13350 = n4103 & n13349;
  assign n13351 = n3740 & n13350;
  assign n13352 = ~n3940 & n13351;
  assign n13353 = ~n4001 & n13352;
  assign n13354 = ~n5043 & n13353;
  assign n13355 = ~n5943 & n13354;
  assign n13356 = ~n6951 & n13355;
  assign n13357 = ~n8037 & n13356;
  assign n13358 = ~n9200 & n13357;
  assign n13359 = ~n13348 & n13358;
  assign n13360 = ~n13347 & n13359;
  assign n13361 = ~n10445 & n13360;
  assign n13362 = ~n12861 & n13361;
  assign n13363 = ~n11846 & n13362;
  assign n13364 = ~n13346 & n13363;
  assign n13365 = n11832 & ~n13076;
  assign n13366 = n11838 & ~n12005;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = n13364 & n13367;
  assign n13369 = n13345 & n13368;
  assign n13370 = n11803 & ~n11928;
  assign n13371 = n11813 & ~n12380;
  assign n13372 = ~n13370 & ~n13371;
  assign n13373 = n11835 & ~n12121;
  assign n13374 = n11834 & ~n12181;
  assign n13375 = ~n13373 & ~n13374;
  assign n13376 = n13372 & n13375;
  assign n13377 = ~n11551 & n11842;
  assign n13378 = n11802 & ~n12158;
  assign n13379 = ~n13377 & ~n13378;
  assign n13380 = ~n11662 & n11839;
  assign n13381 = ~n11588 & n11799;
  assign n13382 = ~n13380 & ~n13381;
  assign n13383 = n13379 & n13382;
  assign n13384 = ~n11611 & n11831;
  assign n13385 = n11812 & ~n12471;
  assign n13386 = ~n13384 & ~n13385;
  assign n13387 = n11811 & ~n13036;
  assign n13388 = n11800 & ~n12240;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = n13386 & n13389;
  assign n13391 = n13383 & n13390;
  assign n13392 = n13376 & n13391;
  assign n13393 = n13369 & n13392;
  assign n13394 = n11847 & ~n13312;
  assign n13395 = ~n13310 & n13394;
  assign n13396 = n13317 & n13395;
  assign n13397 = ~n13393 & ~n13396;
  assign n13398 = ~n13340 & n13397;
  assign n13399 = ~n11662 & n11852;
  assign n13400 = ~n12861 & n12950;
  assign n13401 = ~n13399 & n13400;
  assign n13402 = ~n11846 & n11855;
  assign n13403 = n11857 & ~n13076;
  assign n13404 = n11856 & ~n13036;
  assign n13405 = ~n13403 & ~n13404;
  assign n13406 = ~n13402 & n13405;
  assign n13407 = n13401 & n13406;
  assign n13408 = n3621 & ~n3650;
  assign n13409 = n10462 & n13408;
  assign n13410 = ~n3940 & n13409;
  assign n13411 = ~n4001 & n13410;
  assign n13412 = ~n5043 & n13411;
  assign n13413 = ~n5943 & n13412;
  assign n13414 = ~n6951 & n13413;
  assign n13415 = ~n8037 & n13414;
  assign n13416 = ~n9200 & n13415;
  assign n13417 = ~n13348 & n13416;
  assign n13418 = ~n13347 & n13417;
  assign n13419 = ~n10445 & n13418;
  assign n13420 = ~n12861 & n13419;
  assign n13421 = ~n11846 & n13420;
  assign n13422 = ~n13346 & n13421;
  assign n13423 = n13367 & n13422;
  assign n13424 = n13345 & n13423;
  assign n13425 = n13392 & n13424;
  assign n13426 = ~n13407 & ~n13425;
  assign n13427 = ~n13398 & n13426;
  assign n13428 = ~n11860 & n11881;
  assign n13429 = ~n12861 & n13428;
  assign n13430 = ~n13399 & n13429;
  assign n13431 = n13406 & n13430;
  assign n13432 = n11893 & ~n12041;
  assign n13433 = n11892 & ~n11959;
  assign n13434 = ~n12950 & ~n13433;
  assign n13435 = ~n13432 & n13434;
  assign n13436 = n11897 & ~n12380;
  assign n13437 = n4341 & ~n12902;
  assign n13438 = n4311 & ~n12946;
  assign n13439 = ~n4817 & n10497;
  assign n13440 = ~n4902 & n13439;
  assign n13441 = ~n6001 & n13440;
  assign n13442 = ~n7014 & n13441;
  assign n13443 = ~n8114 & n13442;
  assign n13444 = ~n9276 & n13443;
  assign n13445 = ~n13438 & n13444;
  assign n13446 = ~n13437 & n13445;
  assign n13447 = ~n10523 & n13446;
  assign n13448 = ~n12861 & n13447;
  assign n13449 = ~n11928 & n13448;
  assign n13450 = ~n13436 & n13449;
  assign n13451 = ~n11662 & n11921;
  assign n13452 = n11896 & ~n13076;
  assign n13453 = ~n13451 & ~n13452;
  assign n13454 = n13450 & n13453;
  assign n13455 = n13435 & n13454;
  assign n13456 = n11889 & ~n12158;
  assign n13457 = n11916 & ~n12181;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = ~n11551 & n11914;
  assign n13460 = n11924 & ~n12121;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = n13458 & n13461;
  assign n13463 = n11898 & ~n12471;
  assign n13464 = ~n11588 & n11888;
  assign n13465 = ~n13463 & ~n13464;
  assign n13466 = ~n11846 & n11920;
  assign n13467 = n11923 & ~n12083;
  assign n13468 = ~n13466 & ~n13467;
  assign n13469 = n13465 & n13468;
  assign n13470 = n11886 & ~n12005;
  assign n13471 = ~n11611 & n11917;
  assign n13472 = ~n13470 & ~n13471;
  assign n13473 = n11885 & ~n12240;
  assign n13474 = n11913 & ~n13036;
  assign n13475 = ~n13473 & ~n13474;
  assign n13476 = n13472 & n13475;
  assign n13477 = n13469 & n13476;
  assign n13478 = n13462 & n13477;
  assign n13479 = n13455 & n13478;
  assign n13480 = ~n13431 & ~n13479;
  assign n13481 = ~n13427 & n13480;
  assign n13482 = ~n11928 & n11949;
  assign n13483 = ~n11662 & n11956;
  assign n13484 = n11950 & ~n13076;
  assign n13485 = ~n13483 & ~n13484;
  assign n13486 = ~n13482 & n13485;
  assign n13487 = n12860 & ~n12861;
  assign n13488 = ~n12950 & n13487;
  assign n13489 = n11948 & ~n13036;
  assign n13490 = ~n11846 & n11955;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = n13488 & n13491;
  assign n13493 = n13486 & n13492;
  assign n13494 = ~n4489 & n5084;
  assign n13495 = n10527 & n13494;
  assign n13496 = ~n4817 & n13495;
  assign n13497 = ~n4902 & n13496;
  assign n13498 = ~n6001 & n13497;
  assign n13499 = ~n7014 & n13498;
  assign n13500 = ~n8114 & n13499;
  assign n13501 = ~n9276 & n13500;
  assign n13502 = ~n13438 & n13501;
  assign n13503 = ~n13437 & n13502;
  assign n13504 = ~n10523 & n13503;
  assign n13505 = ~n12861 & n13504;
  assign n13506 = ~n11928 & n13505;
  assign n13507 = ~n13436 & n13506;
  assign n13508 = n13453 & n13507;
  assign n13509 = n13435 & n13508;
  assign n13510 = n13478 & n13509;
  assign n13511 = ~n13493 & ~n13510;
  assign n13512 = ~n13481 & n13511;
  assign n13513 = n11969 & ~n12041;
  assign n13514 = n13094 & ~n13513;
  assign n13515 = n11973 & ~n12380;
  assign n13516 = n5230 & ~n12902;
  assign n13517 = n5598 & ~n12946;
  assign n13518 = n6066 & n6068;
  assign n13519 = ~n5808 & n13518;
  assign n13520 = ~n6056 & n13519;
  assign n13521 = ~n7073 & n13520;
  assign n13522 = ~n8179 & n13521;
  assign n13523 = ~n9344 & n13522;
  assign n13524 = ~n13517 & n13523;
  assign n13525 = ~n13516 & n13524;
  assign n13526 = ~n10594 & n13525;
  assign n13527 = ~n12861 & n13526;
  assign n13528 = ~n12005 & n13527;
  assign n13529 = ~n13515 & n13528;
  assign n13530 = ~n11662 & n11998;
  assign n13531 = n11972 & ~n13076;
  assign n13532 = ~n13530 & ~n13531;
  assign n13533 = n13529 & n13532;
  assign n13534 = n13514 & n13533;
  assign n13535 = n11963 & ~n12158;
  assign n13536 = n11994 & ~n12181;
  assign n13537 = ~n13535 & ~n13536;
  assign n13538 = ~n11551 & n11990;
  assign n13539 = n12001 & ~n12121;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = n13537 & n13540;
  assign n13542 = n11974 & ~n12471;
  assign n13543 = ~n11588 & n11991;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = ~n11846 & n11966;
  assign n13546 = n12000 & ~n12083;
  assign n13547 = ~n13545 & ~n13546;
  assign n13548 = n13544 & n13547;
  assign n13549 = ~n11928 & n11997;
  assign n13550 = ~n11611 & n11993;
  assign n13551 = ~n13549 & ~n13550;
  assign n13552 = n11962 & ~n12240;
  assign n13553 = n11965 & ~n13036;
  assign n13554 = ~n13552 & ~n13553;
  assign n13555 = n13551 & n13554;
  assign n13556 = n13548 & n13555;
  assign n13557 = n13541 & n13556;
  assign n13558 = n13534 & n13557;
  assign n13559 = ~n11959 & n12006;
  assign n13560 = ~n12861 & n13559;
  assign n13561 = ~n12950 & n13560;
  assign n13562 = n13491 & n13561;
  assign n13563 = n13486 & n13562;
  assign n13564 = ~n13558 & ~n13563;
  assign n13565 = ~n13512 & n13564;
  assign n13566 = ~n12005 & n12029;
  assign n13567 = ~n11846 & n12038;
  assign n13568 = ~n13566 & ~n13567;
  assign n13569 = ~n11928 & n12037;
  assign n13570 = ~n11662 & n12028;
  assign n13571 = ~n13569 & ~n13570;
  assign n13572 = n13568 & n13571;
  assign n13573 = ~n12861 & n12951;
  assign n13574 = n13094 & n13573;
  assign n13575 = n12032 & ~n13076;
  assign n13576 = n12031 & ~n13036;
  assign n13577 = ~n13575 & ~n13576;
  assign n13578 = n13574 & n13577;
  assign n13579 = n13572 & n13578;
  assign n13580 = n5379 & ~n5408;
  assign n13581 = ~pi011 & ~n5627;
  assign n13582 = n5687 & n13581;
  assign n13583 = n13580 & n13582;
  assign n13584 = ~n5808 & n13583;
  assign n13585 = ~n6056 & n13584;
  assign n13586 = ~n7073 & n13585;
  assign n13587 = ~n8179 & n13586;
  assign n13588 = ~n9344 & n13587;
  assign n13589 = ~n13517 & n13588;
  assign n13590 = ~n13516 & n13589;
  assign n13591 = ~n10594 & n13590;
  assign n13592 = ~n12861 & n13591;
  assign n13593 = ~n12005 & n13592;
  assign n13594 = ~n13515 & n13593;
  assign n13595 = n13532 & n13594;
  assign n13596 = n13514 & n13595;
  assign n13597 = n13557 & n13596;
  assign n13598 = ~n13579 & ~n13597;
  assign n13599 = ~n13565 & n13598;
  assign n13600 = ~n12005 & n12078;
  assign n13601 = n6672 & ~n12902;
  assign n13602 = n6493 & ~n12946;
  assign n13603 = ~n6522 & ~n6643;
  assign n13604 = n6614 & n13603;
  assign n13605 = n12054 & n13604;
  assign n13606 = ~n6784 & n13605;
  assign n13607 = ~n7158 & n13606;
  assign n13608 = ~n8250 & n13607;
  assign n13609 = ~n9414 & n13608;
  assign n13610 = ~n13602 & n13609;
  assign n13611 = ~n13601 & n13610;
  assign n13612 = ~n10667 & n13611;
  assign n13613 = ~n12861 & n13612;
  assign n13614 = ~n12083 & n13613;
  assign n13615 = ~n13600 & n13614;
  assign n13616 = n12069 & ~n13076;
  assign n13617 = ~n11846 & n12048;
  assign n13618 = ~n13616 & ~n13617;
  assign n13619 = n13615 & n13618;
  assign n13620 = n13095 & n13619;
  assign n13621 = n12045 & ~n12158;
  assign n13622 = n12079 & ~n12121;
  assign n13623 = ~n13621 & ~n13622;
  assign n13624 = n12052 & ~n12380;
  assign n13625 = n12071 & ~n12181;
  assign n13626 = ~n13624 & ~n13625;
  assign n13627 = n13623 & n13626;
  assign n13628 = ~n11551 & n12068;
  assign n13629 = ~n11588 & n12047;
  assign n13630 = ~n13628 & ~n13629;
  assign n13631 = ~n11662 & n12076;
  assign n13632 = n12044 & ~n12240;
  assign n13633 = ~n13631 & ~n13632;
  assign n13634 = n13630 & n13633;
  assign n13635 = ~n11611 & n12072;
  assign n13636 = n12053 & ~n12471;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = n12051 & ~n13036;
  assign n13639 = ~n11928 & n12075;
  assign n13640 = ~n13638 & ~n13639;
  assign n13641 = n13637 & n13640;
  assign n13642 = n13634 & n13641;
  assign n13643 = n13627 & n13642;
  assign n13644 = n13620 & n13643;
  assign n13645 = ~n12041 & n12084;
  assign n13646 = ~n12861 & n13645;
  assign n13647 = n13094 & n13646;
  assign n13648 = n13577 & n13647;
  assign n13649 = n13572 & n13648;
  assign n13650 = ~n13644 & ~n13649;
  assign n13651 = ~n13599 & n13650;
  assign n13652 = n7356 & ~n12946;
  assign n13653 = n7446 & ~n12902;
  assign n13654 = n7752 & n8364;
  assign n13655 = n7693 & n13654;
  assign n13656 = ~n7869 & n13655;
  assign n13657 = ~n8346 & n13656;
  assign n13658 = ~n9485 & n13657;
  assign n13659 = ~n13653 & n13658;
  assign n13660 = ~n13652 & n13659;
  assign n13661 = ~n10741 & n13660;
  assign n13662 = ~n12861 & n13661;
  assign n13663 = ~n12158 & n13662;
  assign n13664 = ~n13052 & n13663;
  assign n13665 = n12130 & ~n12471;
  assign n13666 = ~n11662 & n12153;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = n13664 & n13667;
  assign n13669 = n13095 & n13668;
  assign n13670 = ~n11588 & n12126;
  assign n13671 = n12122 & ~n13036;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = n12147 & ~n12181;
  assign n13674 = ~n11551 & n12144;
  assign n13675 = ~n13673 & ~n13674;
  assign n13676 = n13672 & n13675;
  assign n13677 = ~n11928 & n12151;
  assign n13678 = ~n11611 & n12143;
  assign n13679 = ~n13677 & ~n13678;
  assign n13680 = n12129 & ~n12380;
  assign n13681 = ~n12083 & n12125;
  assign n13682 = ~n13680 & ~n13681;
  assign n13683 = n13679 & n13682;
  assign n13684 = n12123 & ~n12240;
  assign n13685 = ~n11846 & n12150;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = ~n12005 & n12154;
  assign n13688 = n12146 & ~n13076;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = n13686 & n13689;
  assign n13691 = n13683 & n13690;
  assign n13692 = n13676 & n13691;
  assign n13693 = n13669 & n13692;
  assign n13694 = ~n6522 & n7176;
  assign n13695 = n7175 & n10675;
  assign n13696 = n13694 & n13695;
  assign n13697 = ~n6784 & n13696;
  assign n13698 = ~n7158 & n13697;
  assign n13699 = ~n8250 & n13698;
  assign n13700 = ~n9414 & n13699;
  assign n13701 = ~n13602 & n13700;
  assign n13702 = ~n13601 & n13701;
  assign n13703 = ~n10667 & n13702;
  assign n13704 = ~n12861 & n13703;
  assign n13705 = ~n12083 & n13704;
  assign n13706 = ~n13600 & n13705;
  assign n13707 = n13618 & n13706;
  assign n13708 = n13095 & n13707;
  assign n13709 = n13643 & n13708;
  assign n13710 = n12108 & ~n13076;
  assign n13711 = ~n11928 & n12105;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = ~n11662 & n12117;
  assign n13714 = ~n12083 & n12112;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = n13712 & n13715;
  assign n13717 = n12106 & ~n13036;
  assign n13718 = n11501 & ~n12861;
  assign n13719 = ~n12121 & n13718;
  assign n13720 = ~n13717 & n13719;
  assign n13721 = ~n11846 & n12109;
  assign n13722 = ~n12005 & n12116;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = n13720 & n13723;
  assign n13725 = n13095 & n13724;
  assign n13726 = n13716 & n13725;
  assign n13727 = ~n13709 & ~n13726;
  assign n13728 = ~n13693 & n13727;
  assign n13729 = ~n13651 & n13728;
  assign n13730 = ~n7475 & ~n7751;
  assign n13731 = ~n7505 & n13730;
  assign n13732 = n9497 & n13731;
  assign n13733 = ~n7869 & n13732;
  assign n13734 = ~n8346 & n13733;
  assign n13735 = ~n9485 & n13734;
  assign n13736 = ~n13653 & n13735;
  assign n13737 = ~n13652 & n13736;
  assign n13738 = ~n10741 & n13737;
  assign n13739 = ~n12861 & n13738;
  assign n13740 = ~n12158 & n13739;
  assign n13741 = ~n13052 & n13740;
  assign n13742 = n13667 & n13741;
  assign n13743 = n13095 & n13742;
  assign n13744 = n13692 & n13743;
  assign n13745 = ~n11662 & n12165;
  assign n13746 = n12173 & ~n13036;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = ~n12083 & n12162;
  assign n13749 = ~n12158 & n12169;
  assign n13750 = ~n13748 & ~n13749;
  assign n13751 = n13747 & n13750;
  assign n13752 = ~n11928 & n12166;
  assign n13753 = ~n11846 & n12163;
  assign n13754 = ~n13752 & ~n13753;
  assign n13755 = ~n12005 & n12170;
  assign n13756 = n12172 & ~n13076;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = n13754 & n13757;
  assign n13759 = n11478 & ~n12861;
  assign n13760 = ~n12181 & n13759;
  assign n13761 = ~n13052 & n13760;
  assign n13762 = n13095 & n13761;
  assign n13763 = n13758 & n13762;
  assign n13764 = n13751 & n13763;
  assign n13765 = ~n10705 & n12195;
  assign n13766 = ~n12861 & n13765;
  assign n13767 = ~n12121 & n13766;
  assign n13768 = ~n13717 & n13767;
  assign n13769 = n13723 & n13768;
  assign n13770 = n13095 & n13769;
  assign n13771 = n13716 & n13770;
  assign n13772 = ~n13764 & ~n13771;
  assign n13773 = ~n13744 & n13772;
  assign n13774 = ~n13729 & n13773;
  assign n13775 = ~n11318 & n12243;
  assign n13776 = ~n12861 & n13775;
  assign n13777 = ~n12181 & n13776;
  assign n13778 = ~n13052 & n13777;
  assign n13779 = n13095 & n13778;
  assign n13780 = n13758 & n13779;
  assign n13781 = n13751 & n13780;
  assign n13782 = ~n13774 & ~n13781;
  assign n13783 = ~n13135 & ~n13782;
  assign n13784 = ~pi017 & ~n8574;
  assign n13785 = n11377 & n13784;
  assign n13786 = n9942 & n13785;
  assign n13787 = ~n8834 & n13786;
  assign n13788 = ~n10002 & n13787;
  assign n13789 = ~n13097 & n13788;
  assign n13790 = ~n13096 & n13789;
  assign n13791 = ~n11297 & n13790;
  assign n13792 = ~n12861 & n13791;
  assign n13793 = ~n12240 & n13792;
  assign n13794 = ~n12973 & n13793;
  assign n13795 = n13109 & n13794;
  assign n13796 = n13095 & n13795;
  assign n13797 = n13134 & n13796;
  assign n13798 = n11509 & ~n12861;
  assign n13799 = ~n11611 & n13798;
  assign n13800 = ~n12973 & n13799;
  assign n13801 = n11603 & ~n12083;
  assign n13802 = ~n13052 & ~n13801;
  assign n13803 = n13800 & n13802;
  assign n13804 = n13095 & n13803;
  assign n13805 = n11606 & ~n12158;
  assign n13806 = n11599 & ~n13036;
  assign n13807 = ~n13805 & ~n13806;
  assign n13808 = n11596 & ~n12005;
  assign n13809 = n11597 & ~n13076;
  assign n13810 = ~n13808 & ~n13809;
  assign n13811 = n13807 & n13810;
  assign n13812 = n11607 & ~n11928;
  assign n13813 = n11600 & ~n12240;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = n11604 & ~n11662;
  assign n13816 = n11592 & ~n11846;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = n13814 & n13817;
  assign n13819 = n13811 & n13818;
  assign n13820 = n13804 & n13819;
  assign n13821 = ~n13797 & ~n13820;
  assign n13822 = ~n13783 & n13821;
  assign n13823 = n9622 & ~n12946;
  assign n13824 = n9687 & ~n12902;
  assign n13825 = ~n9717 & ~n9913;
  assign n13826 = n9856 & n13825;
  assign n13827 = ~n9929 & n13826;
  assign n13828 = ~n13824 & n13827;
  assign n13829 = ~n13823 & n13828;
  assign n13830 = ~n11266 & n13829;
  assign n13831 = ~n12861 & n13830;
  assign n13832 = ~n11588 & n13831;
  assign n13833 = ~n12973 & n13832;
  assign n13834 = n13054 & n13833;
  assign n13835 = n13095 & n13834;
  assign n13836 = n11580 & ~n12083;
  assign n13837 = n11583 & ~n12240;
  assign n13838 = ~n13836 & ~n13837;
  assign n13839 = n11577 & ~n11662;
  assign n13840 = n11576 & ~n12158;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = n13838 & n13841;
  assign n13843 = n11584 & ~n12005;
  assign n13844 = n11554 & ~n13076;
  assign n13845 = ~n13843 & ~n13844;
  assign n13846 = n11581 & ~n11928;
  assign n13847 = n11553 & ~n11846;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = n13845 & n13848;
  assign n13850 = n11557 & ~n12380;
  assign n13851 = ~n11551 & n11574;
  assign n13852 = ~n13850 & ~n13851;
  assign n13853 = n11573 & ~n13036;
  assign n13854 = n11558 & ~n12471;
  assign n13855 = ~n13853 & ~n13854;
  assign n13856 = n13852 & n13855;
  assign n13857 = n13849 & n13856;
  assign n13858 = n13842 & n13857;
  assign n13859 = n13835 & n13858;
  assign n13860 = ~n10787 & n12266;
  assign n13861 = ~n12861 & n13860;
  assign n13862 = ~n11611 & n13861;
  assign n13863 = ~n12973 & n13862;
  assign n13864 = n13802 & n13863;
  assign n13865 = n13095 & n13864;
  assign n13866 = n13819 & n13865;
  assign n13867 = ~n13859 & ~n13866;
  assign n13868 = ~n13822 & n13867;
  assign n13869 = ~pi019 & ~n9717;
  assign n13870 = ~n9913 & n13869;
  assign n13871 = n9856 & n13870;
  assign n13872 = ~n9929 & n13871;
  assign n13873 = ~n13824 & n13872;
  assign n13874 = ~n13823 & n13873;
  assign n13875 = ~n11266 & n13874;
  assign n13876 = ~n12861 & n13875;
  assign n13877 = ~n11588 & n13876;
  assign n13878 = ~n12973 & n13877;
  assign n13879 = n13054 & n13878;
  assign n13880 = n13095 & n13879;
  assign n13881 = n13858 & n13880;
  assign n13882 = n11479 & ~n11588;
  assign n13883 = n11537 & ~n13036;
  assign n13884 = ~n13882 & ~n13883;
  assign n13885 = n13054 & n13884;
  assign n13886 = n12376 & ~n12861;
  assign n13887 = ~n11551 & n13886;
  assign n13888 = ~n12973 & n13887;
  assign n13889 = n13095 & n13888;
  assign n13890 = n13885 & n13889;
  assign n13891 = n11516 & ~n12158;
  assign n13892 = n11540 & ~n12240;
  assign n13893 = ~n13891 & ~n13892;
  assign n13894 = n11500 & ~n13076;
  assign n13895 = n11543 & ~n11928;
  assign n13896 = ~n13894 & ~n13895;
  assign n13897 = n13893 & n13896;
  assign n13898 = n11544 & ~n11662;
  assign n13899 = n11539 & ~n12083;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = n11547 & ~n12005;
  assign n13902 = n11546 & ~n11846;
  assign n13903 = ~n13901 & ~n13902;
  assign n13904 = n13900 & n13903;
  assign n13905 = n13897 & n13904;
  assign n13906 = n13890 & n13905;
  assign n13907 = ~n13881 & ~n13906;
  assign n13908 = n12641 & ~n12946;
  assign n13909 = ~n12671 & ~n12811;
  assign n13910 = ~n12743 & ~n12841;
  assign n13911 = ~n12713 & ~n12773;
  assign n13912 = n13910 & n13911;
  assign n13913 = n13909 & n13912;
  assign n13914 = ~n12902 & n13913;
  assign n13915 = ~n13908 & n13914;
  assign n13916 = ~n12861 & n13915;
  assign n13917 = ~n12860 & n13916;
  assign n13918 = n12952 & n13917;
  assign n13919 = n12974 & n13054;
  assign n13920 = n13918 & n13919;
  assign n13921 = ~n2754 & ~n3066;
  assign n13922 = ~n3983 & n13921;
  assign n13923 = ~n4024 & n13922;
  assign n13924 = ~n4999 & n13923;
  assign n13925 = ~n5827 & n13924;
  assign n13926 = ~n6893 & n13925;
  assign n13927 = ~n7890 & n13926;
  assign n13928 = ~n9131 & n13927;
  assign n13929 = ~n10278 & n13928;
  assign n13930 = ~n11662 & n13929;
  assign n13931 = ~n9687 & ~n9929;
  assign n13932 = ~n11266 & n13931;
  assign n13933 = ~n11588 & n13932;
  assign n13934 = ~n13930 & ~n13933;
  assign n13935 = ~n4341 & ~n4817;
  assign n13936 = ~n4902 & n13935;
  assign n13937 = ~n6001 & n13936;
  assign n13938 = ~n7014 & n13937;
  assign n13939 = ~n8114 & n13938;
  assign n13940 = ~n9276 & n13939;
  assign n13941 = ~n10523 & n13940;
  assign n13942 = ~n11928 & n13941;
  assign n13943 = ~n5230 & ~n5808;
  assign n13944 = ~n6056 & n13943;
  assign n13945 = ~n7073 & n13944;
  assign n13946 = ~n8179 & n13945;
  assign n13947 = ~n9344 & n13946;
  assign n13948 = ~n10594 & n13947;
  assign n13949 = ~n12005 & n13948;
  assign n13950 = ~n13942 & ~n13949;
  assign n13951 = n13934 & n13950;
  assign n13952 = ~n841 & ~n1372;
  assign n13953 = ~n2243 & n13952;
  assign n13954 = ~n3104 & n13953;
  assign n13955 = ~n3971 & n13954;
  assign n13956 = ~n4872 & n13955;
  assign n13957 = ~n5801 & n13956;
  assign n13958 = ~n6739 & n13957;
  assign n13959 = ~n7807 & n13958;
  assign n13960 = ~n8989 & n13959;
  assign n13961 = ~n10273 & n13960;
  assign n13962 = ~n11499 & n13961;
  assign n13963 = ~n13076 & n13962;
  assign n13964 = ~n3798 & ~n3940;
  assign n13965 = ~n4001 & n13964;
  assign n13966 = ~n5043 & n13965;
  assign n13967 = ~n5943 & n13966;
  assign n13968 = ~n6951 & n13967;
  assign n13969 = ~n8037 & n13968;
  assign n13970 = ~n9200 & n13969;
  assign n13971 = ~n10445 & n13970;
  assign n13972 = ~n11846 & n13971;
  assign n13973 = ~n13963 & ~n13972;
  assign n13974 = ~n7446 & ~n7869;
  assign n13975 = ~n8346 & n13974;
  assign n13976 = ~n9485 & n13975;
  assign n13977 = ~n10741 & n13976;
  assign n13978 = ~n12158 & n13977;
  assign n13979 = ~n8603 & ~n8834;
  assign n13980 = ~n10002 & n13979;
  assign n13981 = ~n11297 & n13980;
  assign n13982 = ~n12240 & n13981;
  assign n13983 = ~n13978 & ~n13982;
  assign n13984 = n13973 & n13983;
  assign n13985 = ~n6672 & ~n6784;
  assign n13986 = ~n7158 & n13985;
  assign n13987 = ~n8250 & n13986;
  assign n13988 = ~n9414 & n13987;
  assign n13989 = ~n10667 & n13988;
  assign n13990 = ~n12083 & n13989;
  assign n13991 = ~n13055 & ~n13990;
  assign n13992 = ~n1617 & ~n2242;
  assign n13993 = ~n3095 & n13992;
  assign n13994 = ~n3997 & n13993;
  assign n13995 = ~n4837 & n13994;
  assign n13996 = ~n5822 & n13995;
  assign n13997 = ~n6820 & n13996;
  assign n13998 = ~n7785 & n13997;
  assign n13999 = ~n9027 & n13998;
  assign n14000 = ~n10245 & n13999;
  assign n14001 = ~n11536 & n14000;
  assign n14002 = ~n13036 & n14001;
  assign n14003 = ~n10939 & ~n11188;
  assign n14004 = ~n12380 & n14003;
  assign n14005 = ~n14002 & ~n14004;
  assign n14006 = n13991 & n14005;
  assign n14007 = n13984 & n14006;
  assign n14008 = n13951 & n14007;
  assign n14009 = n13920 & n14008;
  assign n14010 = n10969 & ~n12946;
  assign n14011 = n10939 & ~n12902;
  assign n14012 = ~n10909 & ~n11168;
  assign n14013 = n11135 & n14012;
  assign n14014 = ~n11188 & n14013;
  assign n14015 = ~n14011 & n14014;
  assign n14016 = ~n14010 & n14015;
  assign n14017 = ~n12861 & n14016;
  assign n14018 = ~n12380 & n14017;
  assign n14019 = ~n12972 & n14018;
  assign n14020 = ~n12973 & ~n13052;
  assign n14021 = n14019 & n14020;
  assign n14022 = n13095 & n14021;
  assign n14023 = ~n12240 & n12311;
  assign n14024 = ~n11928 & n12308;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = ~n11846 & n12335;
  assign n14027 = ~n12005 & n12364;
  assign n14028 = ~n14026 & ~n14027;
  assign n14029 = n14025 & n14028;
  assign n14030 = ~n12158 & n12347;
  assign n14031 = ~n12083 & n12340;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = n12375 & ~n13036;
  assign n14034 = n12300 & ~n13076;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = n14032 & n14035;
  assign n14037 = n12314 & ~n12471;
  assign n14038 = ~n13053 & ~n14037;
  assign n14039 = ~n11588 & n12343;
  assign n14040 = ~n11662 & n12358;
  assign n14041 = ~n14039 & ~n14040;
  assign n14042 = n14038 & n14041;
  assign n14043 = n14036 & n14042;
  assign n14044 = n14029 & n14043;
  assign n14045 = n14022 & n14044;
  assign n14046 = ~n10879 & ~n12861;
  assign n14047 = ~n12471 & n14046;
  assign n14048 = ~n12972 & n14047;
  assign n14049 = n14020 & n14048;
  assign n14050 = n13095 & n14049;
  assign n14051 = ~n12083 & n12461;
  assign n14052 = n12401 & ~n13076;
  assign n14053 = ~n14051 & ~n14052;
  assign n14054 = ~n11846 & n12409;
  assign n14055 = ~n12380 & n12412;
  assign n14056 = ~n14054 & ~n14055;
  assign n14057 = n14053 & n14056;
  assign n14058 = ~n12158 & n12466;
  assign n14059 = ~n12005 & n12435;
  assign n14060 = ~n14058 & ~n14059;
  assign n14061 = n12456 & ~n13036;
  assign n14062 = ~n11588 & n12467;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = n14060 & n14063;
  assign n14065 = ~n11662 & n12444;
  assign n14066 = ~n13053 & ~n14065;
  assign n14067 = ~n12240 & n12421;
  assign n14068 = ~n11928 & n12428;
  assign n14069 = ~n14067 & ~n14068;
  assign n14070 = n14066 & n14069;
  assign n14071 = n14064 & n14070;
  assign n14072 = n14057 & n14071;
  assign n14073 = n14050 & n14072;
  assign n14074 = ~n14045 & ~n14073;
  assign n14075 = ~n14009 & n14074;
  assign n14076 = n13907 & n14075;
  assign n14077 = ~n13868 & n14076;
  assign n14078 = n12487 & ~n12861;
  assign n14079 = ~n12471 & n14078;
  assign n14080 = ~n12972 & n14079;
  assign n14081 = n14020 & n14080;
  assign n14082 = n13095 & n14081;
  assign n14083 = n14072 & n14082;
  assign n14084 = ~n11343 & n12381;
  assign n14085 = ~n12861 & n14084;
  assign n14086 = ~n11551 & n14085;
  assign n14087 = ~n12973 & n14086;
  assign n14088 = n13095 & n14087;
  assign n14089 = n13885 & n14088;
  assign n14090 = n13905 & n14089;
  assign n14091 = ~n14083 & ~n14090;
  assign n14092 = pi021 & ~n10909;
  assign n14093 = ~n11168 & n14092;
  assign n14094 = n11135 & n14093;
  assign n14095 = ~n11188 & n14094;
  assign n14096 = ~n14011 & n14095;
  assign n14097 = ~n14010 & n14096;
  assign n14098 = ~n12861 & n14097;
  assign n14099 = ~n12380 & n14098;
  assign n14100 = ~n12972 & n14099;
  assign n14101 = n14020 & n14100;
  assign n14102 = n13095 & n14101;
  assign n14103 = n14044 & n14102;
  assign n14104 = pi023 & ~n12671;
  assign n14105 = ~n12811 & n14104;
  assign n14106 = n13912 & n14105;
  assign n14107 = ~n12902 & n14106;
  assign n14108 = ~n13908 & n14107;
  assign n14109 = ~n12861 & n14108;
  assign n14110 = ~n12860 & n14109;
  assign n14111 = n12952 & n14110;
  assign n14112 = n13919 & n14111;
  assign n14113 = n14008 & n14112;
  assign n14114 = ~n14103 & ~n14113;
  assign n14115 = n14091 & n14114;
  assign n14116 = ~n14077 & n14115;
  assign n14117 = ~n13093 & ~n14116;
  assign n14118 = pi024 & ~n12946;
  assign n14119 = ~n12903 & n14118;
  assign n14120 = ~n12861 & n14119;
  assign n14121 = ~n12860 & n14120;
  assign n14122 = n12952 & n14121;
  assign n14123 = n12975 & n14122;
  assign n14124 = n13092 & n14123;
  assign n14125 = ~n7223 & ~n7295;
  assign n14126 = ~n7218 & ~n7229;
  assign n14127 = n14125 & n14126;
  assign n14128 = ~n6492 & ~n6521;
  assign n14129 = n10826 & n14128;
  assign n14130 = n6182 & n14129;
  assign n14131 = ~n8542 & n12537;
  assign n14132 = ~n7355 & ~n7750;
  assign n14133 = n10824 & n14132;
  assign n14134 = n14131 & n14133;
  assign n14135 = n14130 & n14134;
  assign n14136 = ~n3372 & ~n3738;
  assign n14137 = ~n3283 & ~n3402;
  assign n14138 = n14136 & n14137;
  assign n14139 = n10858 & n12571;
  assign n14140 = n14138 & n14139;
  assign n14141 = ~n4310 & ~n4706;
  assign n14142 = n10828 & n14141;
  assign n14143 = ~n2423 & ~n3254;
  assign n14144 = ~n5377 & ~n5597;
  assign n14145 = n14143 & n14144;
  assign n14146 = n14142 & n14145;
  assign n14147 = n14140 & n14146;
  assign n14148 = n14135 & n14147;
  assign n14149 = ~pi233 & pi241;
  assign n14150 = pi233 & ~pi241;
  assign n14151 = ~pi234 & pi242;
  assign n14152 = pi234 & ~pi242;
  assign n14153 = ~pi235 & pi243;
  assign n14154 = pi235 & ~pi243;
  assign n14155 = ~pi236 & pi244;
  assign n14156 = pi236 & ~pi244;
  assign n14157 = pi238 & ~pi246;
  assign n14158 = pi237 & ~pi245;
  assign n14159 = ~n14157 & ~n14158;
  assign n14160 = ~pi237 & pi245;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n14156 & ~n14161;
  assign n14163 = ~n14155 & ~n14162;
  assign n14164 = ~n14154 & ~n14163;
  assign n14165 = ~n14153 & ~n14164;
  assign n14166 = ~n14152 & ~n14165;
  assign n14167 = ~n14151 & ~n14166;
  assign n14168 = ~n14150 & ~n14167;
  assign n14169 = ~n14149 & ~n14168;
  assign n14170 = ~pi232 & ~n14169;
  assign n14171 = ~pi240 & ~n14170;
  assign n14172 = pi231 & ~pi239;
  assign n14173 = pi232 & ~n14149;
  assign n14174 = ~n14168 & n14173;
  assign n14175 = ~n14172 & ~n14174;
  assign n14176 = ~n14171 & n14175;
  assign n14177 = n12811 & ~n14176;
  assign n14178 = n9824 & n11133;
  assign n14179 = n14177 & n14178;
  assign n14180 = n14148 & n14179;
  assign n14181 = ~n1678 & ~n9651;
  assign n14182 = n12496 & n14181;
  assign n14183 = n12534 & n14182;
  assign n14184 = n12531 & n14183;
  assign n14185 = ~n562 & ~n687;
  assign n14186 = n12582 & n14185;
  assign n14187 = pi026 & ~n501;
  assign n14188 = n12554 & n12872;
  assign n14189 = n14187 & n14188;
  assign n14190 = n11409 & n12916;
  assign n14191 = ~n566 & ~n659;
  assign n14192 = n4792 & n14191;
  assign n14193 = n14190 & n14192;
  assign n14194 = ~n2396 & ~n2484;
  assign n14195 = n12549 & n14194;
  assign n14196 = ~n1404 & ~n1650;
  assign n14197 = n2308 & n14196;
  assign n14198 = n14195 & n14197;
  assign n14199 = n14193 & n14198;
  assign n14200 = n14189 & n14199;
  assign n14201 = ~n6494 & ~n7723;
  assign n14202 = n12544 & n14201;
  assign n14203 = n7242 & n14202;
  assign n14204 = ~pi231 & pi239;
  assign n14205 = ~n8515 & ~n8734;
  assign n14206 = ~n14204 & n14205;
  assign n14207 = n11400 & n12545;
  assign n14208 = n14206 & n14207;
  assign n14209 = n14203 & n14208;
  assign n14210 = ~n2664 & ~n3345;
  assign n14211 = ~n3285 & ~n3711;
  assign n14212 = n14210 & n14211;
  assign n14213 = n6142 & n14212;
  assign n14214 = ~n4679 & ~n5350;
  assign n14215 = n12550 & n14214;
  assign n14216 = n11402 & n14215;
  assign n14217 = n14213 & n14216;
  assign n14218 = n14209 & n14217;
  assign n14219 = n14200 & n14218;
  assign n14220 = ~n1172 & n14219;
  assign n14221 = ~n996 & n14220;
  assign n14222 = ~n2306 & n14221;
  assign n14223 = n3819 & n14222;
  assign n14224 = n3821 & n14223;
  assign n14225 = n14186 & n14224;
  assign n14226 = ~n1432 & ~n1463;
  assign n14227 = n10820 & n14226;
  assign n14228 = n2222 & n12498;
  assign n14229 = n14227 & n14228;
  assign n14230 = n14225 & n14229;
  assign n14231 = n14184 & n14230;
  assign n14232 = n14180 & n14231;
  assign n14233 = ~n7236 & n14232;
  assign n14234 = ~n6137 & n14233;
  assign n14235 = n6193 & n14234;
  assign n14236 = n6134 & n14235;
  assign n14237 = ~n8867 & n14236;
  assign n14238 = ~n8513 & n12537;
  assign n14239 = ~n6612 & ~n7721;
  assign n14240 = n10824 & n14239;
  assign n14241 = n12540 & n14240;
  assign n14242 = n14238 & n14241;
  assign n14243 = ~n2630 & ~n3254;
  assign n14244 = ~n5407 & ~n5597;
  assign n14245 = n14243 & n14244;
  assign n14246 = ~n3372 & ~n3768;
  assign n14247 = n14137 & n14246;
  assign n14248 = n14245 & n14247;
  assign n14249 = ~n4310 & ~n4735;
  assign n14250 = n10828 & n14249;
  assign n14251 = n6182 & n14250;
  assign n14252 = n14248 & n14251;
  assign n14253 = n4792 & n12554;
  assign n14254 = pi025 & ~n501;
  assign n14255 = ~n566 & ~n689;
  assign n14256 = n14254 & n14255;
  assign n14257 = n14253 & n14256;
  assign n14258 = ~n1404 & ~n1681;
  assign n14259 = n12916 & n14258;
  assign n14260 = n12873 & n14259;
  assign n14261 = ~n2484 & ~n2603;
  assign n14262 = ~n3285 & ~n3741;
  assign n14263 = n14261 & n14262;
  assign n14264 = n5716 & n14263;
  assign n14265 = n14260 & n14264;
  assign n14266 = n14257 & n14265;
  assign n14267 = ~n8486 & ~n8734;
  assign n14268 = n11400 & n14267;
  assign n14269 = ~n7328 & ~n7694;
  assign n14270 = n11399 & n14269;
  assign n14271 = ~n6465 & ~n6585;
  assign n14272 = n7241 & n14271;
  assign n14273 = n14270 & n14272;
  assign n14274 = n14268 & n14273;
  assign n14275 = n5722 & n14210;
  assign n14276 = n5721 & n14275;
  assign n14277 = ~n4708 & ~n5380;
  assign n14278 = n10836 & n14277;
  assign n14279 = n12551 & n14278;
  assign n14280 = n14276 & n14279;
  assign n14281 = n14274 & n14280;
  assign n14282 = n14266 & n14281;
  assign n14283 = ~n1172 & n14282;
  assign n14284 = ~n996 & n14283;
  assign n14285 = ~n2306 & n14284;
  assign n14286 = n3819 & n14285;
  assign n14287 = n14139 & n14286;
  assign n14288 = n12583 & n14287;
  assign n14289 = n14252 & n14288;
  assign n14290 = n14242 & n14289;
  assign n14291 = ~pi231 & pi247;
  assign n14292 = ~pi233 & pi249;
  assign n14293 = pi233 & ~pi249;
  assign n14294 = ~pi234 & pi250;
  assign n14295 = pi234 & ~pi250;
  assign n14296 = ~pi235 & pi251;
  assign n14297 = pi235 & ~pi251;
  assign n14298 = ~pi236 & pi252;
  assign n14299 = pi236 & ~pi252;
  assign n14300 = pi238 & ~pi254;
  assign n14301 = pi237 & ~pi253;
  assign n14302 = ~n14300 & ~n14301;
  assign n14303 = ~pi237 & pi253;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = ~n14299 & ~n14304;
  assign n14306 = ~n14298 & ~n14305;
  assign n14307 = ~n14297 & ~n14306;
  assign n14308 = ~n14296 & ~n14307;
  assign n14309 = ~n14295 & ~n14308;
  assign n14310 = ~n14294 & ~n14309;
  assign n14311 = ~n14293 & ~n14310;
  assign n14312 = ~n14292 & ~n14311;
  assign n14313 = ~pi232 & ~n14312;
  assign n14314 = ~pi248 & ~n14313;
  assign n14315 = pi231 & ~pi247;
  assign n14316 = pi232 & ~n14292;
  assign n14317 = ~n14311 & n14316;
  assign n14318 = ~n14315 & ~n14317;
  assign n14319 = ~n14314 & n14318;
  assign n14320 = ~n14291 & ~n14319;
  assign n14321 = ~pi231 & pi271;
  assign n14322 = ~pi233 & pi273;
  assign n14323 = pi233 & ~pi273;
  assign n14324 = ~pi234 & pi274;
  assign n14325 = pi234 & ~pi274;
  assign n14326 = ~pi235 & pi275;
  assign n14327 = pi235 & ~pi275;
  assign n14328 = ~pi236 & pi276;
  assign n14329 = pi236 & ~pi276;
  assign n14330 = pi238 & ~pi278;
  assign n14331 = pi237 & ~pi277;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = ~pi237 & pi277;
  assign n14334 = ~n14332 & ~n14333;
  assign n14335 = ~n14329 & ~n14334;
  assign n14336 = ~n14328 & ~n14335;
  assign n14337 = ~n14327 & ~n14336;
  assign n14338 = ~n14326 & ~n14337;
  assign n14339 = ~n14325 & ~n14338;
  assign n14340 = ~n14324 & ~n14339;
  assign n14341 = ~n14323 & ~n14340;
  assign n14342 = ~n14322 & ~n14341;
  assign n14343 = ~pi232 & ~n14342;
  assign n14344 = ~pi272 & ~n14343;
  assign n14345 = pi231 & ~pi271;
  assign n14346 = pi232 & ~n14322;
  assign n14347 = ~n14341 & n14346;
  assign n14348 = ~n14345 & ~n14347;
  assign n14349 = ~n14344 & n14348;
  assign n14350 = ~n14321 & ~n14349;
  assign n14351 = ~n14320 & ~n14350;
  assign n14352 = ~pi231 & pi263;
  assign n14353 = ~pi233 & pi265;
  assign n14354 = pi233 & ~pi265;
  assign n14355 = ~pi234 & pi266;
  assign n14356 = pi234 & ~pi266;
  assign n14357 = ~pi235 & pi267;
  assign n14358 = pi235 & ~pi267;
  assign n14359 = ~pi236 & pi268;
  assign n14360 = pi236 & ~pi268;
  assign n14361 = pi238 & ~pi270;
  assign n14362 = pi237 & ~pi269;
  assign n14363 = ~n14361 & ~n14362;
  assign n14364 = ~pi237 & pi269;
  assign n14365 = ~n14363 & ~n14364;
  assign n14366 = ~n14360 & ~n14365;
  assign n14367 = ~n14359 & ~n14366;
  assign n14368 = ~n14358 & ~n14367;
  assign n14369 = ~n14357 & ~n14368;
  assign n14370 = ~n14356 & ~n14369;
  assign n14371 = ~n14355 & ~n14370;
  assign n14372 = ~n14354 & ~n14371;
  assign n14373 = ~n14353 & ~n14372;
  assign n14374 = ~pi232 & ~n14373;
  assign n14375 = ~pi264 & ~n14374;
  assign n14376 = pi231 & ~pi263;
  assign n14377 = pi232 & ~n14353;
  assign n14378 = ~n14372 & n14377;
  assign n14379 = ~n14376 & ~n14378;
  assign n14380 = ~n14375 & n14379;
  assign n14381 = ~n14352 & ~n14380;
  assign n14382 = ~n14176 & ~n14204;
  assign n14383 = ~n14381 & ~n14382;
  assign n14384 = n14351 & n14383;
  assign n14385 = n10909 & n12530;
  assign n14386 = n12534 & n14385;
  assign n14387 = ~pi231 & pi255;
  assign n14388 = ~pi233 & pi257;
  assign n14389 = pi233 & ~pi257;
  assign n14390 = ~pi234 & pi258;
  assign n14391 = pi234 & ~pi258;
  assign n14392 = ~pi235 & pi259;
  assign n14393 = pi235 & ~pi259;
  assign n14394 = ~pi236 & pi260;
  assign n14395 = pi236 & ~pi260;
  assign n14396 = pi238 & ~pi262;
  assign n14397 = pi237 & ~pi261;
  assign n14398 = ~n14396 & ~n14397;
  assign n14399 = ~pi237 & pi261;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = ~n14395 & ~n14400;
  assign n14402 = ~n14394 & ~n14401;
  assign n14403 = ~n14393 & ~n14402;
  assign n14404 = ~n14392 & ~n14403;
  assign n14405 = ~n14391 & ~n14404;
  assign n14406 = ~n14390 & ~n14405;
  assign n14407 = ~n14389 & ~n14406;
  assign n14408 = ~n14388 & ~n14407;
  assign n14409 = ~pi232 & ~n14408;
  assign n14410 = ~pi256 & ~n14409;
  assign n14411 = pi231 & ~pi255;
  assign n14412 = pi232 & ~n14388;
  assign n14413 = ~n14407 & n14412;
  assign n14414 = ~n14411 & ~n14413;
  assign n14415 = ~n14410 & n14414;
  assign n14416 = ~n14387 & ~n14415;
  assign n14417 = ~n12526 & ~n12668;
  assign n14418 = ~n12670 & n14417;
  assign n14419 = ~n14416 & n14418;
  assign n14420 = n14386 & n14419;
  assign n14421 = n10820 & n12498;
  assign n14422 = ~n562 & ~n717;
  assign n14423 = n2222 & n14422;
  assign n14424 = n14421 & n14423;
  assign n14425 = n9717 & n12496;
  assign n14426 = ~n1709 & ~n9651;
  assign n14427 = n14226 & n14426;
  assign n14428 = n14425 & n14427;
  assign n14429 = n14424 & n14428;
  assign n14430 = n14420 & n14429;
  assign n14431 = n14384 & n14430;
  assign n14432 = n14290 & n14431;
  assign n14433 = ~n7236 & n14432;
  assign n14434 = ~n6137 & n14433;
  assign n14435 = n6193 & n14434;
  assign n14436 = n6134 & n14435;
  assign n14437 = ~n8867 & n14436;
  assign n14438 = ~n14237 & ~n14437;
  assign n14439 = n11466 & ~n14438;
  assign n14440 = n14127 & n14439;
  assign n14441 = ~n10027 & n14440;
  assign n14442 = ~n8866 & n14441;
  assign n14443 = n8898 & n14442;
  assign n14444 = n8863 & n14443;
  assign n14445 = ~n10788 & n14444;
  assign n14446 = ~n10026 & n14445;
  assign n14447 = n10072 & n14446;
  assign n14448 = n10021 & n14447;
  assign n14449 = ~n14124 & ~n14448;
  assign po013 = n14117 | ~n14449;
  assign n14451 = n12972 & ~n13906;
  assign n14452 = n13053 & ~n13820;
  assign n14453 = ~n14451 & ~n14452;
  assign n14454 = n12973 & ~n13764;
  assign n14455 = n13052 & ~n13726;
  assign n14456 = ~n14454 & ~n14455;
  assign n14457 = n14453 & n14456;
  assign n14458 = ~n5378 & ~n5808;
  assign n14459 = ~n6056 & n14458;
  assign n14460 = ~n7073 & n14459;
  assign n14461 = ~n8179 & n14460;
  assign n14462 = ~n9344 & n14461;
  assign n14463 = ~n10594 & n14462;
  assign n14464 = ~n12005 & n14463;
  assign n14465 = ~n13558 & n14464;
  assign n14466 = n12951 & ~n13579;
  assign n14467 = n12861 & ~n13318;
  assign n14468 = ~n689 & ~n969;
  assign n14469 = n2246 & n14468;
  assign n14470 = n12555 & n14469;
  assign n14471 = ~n1435 & ~n1681;
  assign n14472 = n12559 & n14471;
  assign n14473 = n10841 & n12562;
  assign n14474 = n14472 & n14473;
  assign n14475 = n10845 & n14210;
  assign n14476 = n3942 & n14475;
  assign n14477 = n14474 & n14476;
  assign n14478 = n14470 & n14477;
  assign n14479 = ~n8486 & n12904;
  assign n14480 = n10832 & n14269;
  assign n14481 = ~n6585 & ~n7240;
  assign n14482 = n12544 & n14481;
  assign n14483 = n14480 & n14482;
  assign n14484 = n14479 & n14483;
  assign n14485 = ~n2603 & ~n3227;
  assign n14486 = n12550 & n14485;
  assign n14487 = ~n2635 & ~n3741;
  assign n14488 = ~n3256 & ~n3375;
  assign n14489 = n14487 & n14488;
  assign n14490 = n14486 & n14489;
  assign n14491 = n6741 & n14278;
  assign n14492 = n14490 & n14491;
  assign n14493 = n14484 & n14492;
  assign n14494 = n14478 & n14493;
  assign n14495 = ~n1172 & n14494;
  assign n14496 = ~n996 & n14495;
  assign n14497 = ~n2306 & n14496;
  assign n14498 = n3819 & n14497;
  assign n14499 = n14139 & n14498;
  assign n14500 = n12583 & n14499;
  assign n14501 = n14252 & n14500;
  assign n14502 = n14242 & n14501;
  assign n14503 = n14431 & n14502;
  assign n14504 = ~n7236 & n14503;
  assign n14505 = ~n6137 & n14504;
  assign n14506 = n6193 & n14505;
  assign n14507 = n6134 & n14506;
  assign n14508 = ~n8867 & n14507;
  assign n14509 = ~n7235 & n14508;
  assign n14510 = n7296 & n14509;
  assign n14511 = n7231 & n14510;
  assign n14512 = ~n10027 & n14511;
  assign n14513 = ~n8866 & n14512;
  assign n14514 = n8898 & n14513;
  assign n14515 = n8863 & n14514;
  assign n14516 = ~n10788 & n14515;
  assign n14517 = ~n10026 & n14516;
  assign n14518 = n10072 & n14517;
  assign n14519 = n10021 & n14518;
  assign n14520 = ~n14382 & ~n14519;
  assign n14521 = ~n659 & ~n969;
  assign n14522 = n2246 & n14521;
  assign n14523 = n12555 & n14522;
  assign n14524 = ~n1435 & ~n1650;
  assign n14525 = n12559 & n14524;
  assign n14526 = n14473 & n14525;
  assign n14527 = n14476 & n14526;
  assign n14528 = n14523 & n14527;
  assign n14529 = ~n8515 & ~n14204;
  assign n14530 = n12904 & n14529;
  assign n14531 = n8868 & n14201;
  assign n14532 = n12546 & n14531;
  assign n14533 = n14530 & n14532;
  assign n14534 = ~n2396 & ~n3227;
  assign n14535 = n12550 & n14534;
  assign n14536 = ~n2635 & ~n3711;
  assign n14537 = n14488 & n14536;
  assign n14538 = n14535 & n14537;
  assign n14539 = n10836 & n14214;
  assign n14540 = n6741 & n14539;
  assign n14541 = n14538 & n14540;
  assign n14542 = n14533 & n14541;
  assign n14543 = n14528 & n14542;
  assign n14544 = ~n1172 & n14543;
  assign n14545 = ~n996 & n14544;
  assign n14546 = ~n2306 & n14545;
  assign n14547 = n3819 & n14546;
  assign n14548 = n3821 & n14547;
  assign n14549 = n14186 & n14548;
  assign n14550 = n14229 & n14549;
  assign n14551 = n14184 & n14550;
  assign n14552 = n14180 & n14551;
  assign n14553 = ~n7236 & n14552;
  assign n14554 = ~n6137 & n14553;
  assign n14555 = n6193 & n14554;
  assign n14556 = n6134 & n14555;
  assign n14557 = ~n8867 & n14556;
  assign n14558 = ~n7235 & n14557;
  assign n14559 = n7296 & n14558;
  assign n14560 = n7231 & n14559;
  assign n14561 = ~n10027 & n14560;
  assign n14562 = ~n8866 & n14561;
  assign n14563 = n8898 & n14562;
  assign n14564 = n8863 & n14563;
  assign n14565 = ~n10788 & n14564;
  assign n14566 = ~n10026 & n14565;
  assign n14567 = n10072 & n14566;
  assign n14568 = n10021 & n14567;
  assign n14569 = ~n14520 & ~n14568;
  assign n14570 = ~n14467 & n14569;
  assign n14571 = ~n14466 & n14570;
  assign n14572 = n12860 & ~n13493;
  assign n14573 = n12950 & ~n13407;
  assign n14574 = ~n14572 & ~n14573;
  assign n14575 = n14571 & n14574;
  assign n14576 = ~n14465 & n14575;
  assign n14577 = n13055 & ~n14073;
  assign n14578 = ~n11133 & ~n11188;
  assign n14579 = ~n12380 & n14578;
  assign n14580 = ~n14045 & n14579;
  assign n14581 = ~n14577 & ~n14580;
  assign n14582 = n14576 & n14581;
  assign n14583 = n14457 & n14582;
  assign n14584 = ~n4707 & ~n4817;
  assign n14585 = ~n4902 & n14584;
  assign n14586 = ~n6001 & n14585;
  assign n14587 = ~n7014 & n14586;
  assign n14588 = ~n8114 & n14587;
  assign n14589 = ~n9276 & n14588;
  assign n14590 = ~n10523 & n14589;
  assign n14591 = ~n11928 & n14590;
  assign n14592 = ~n13479 & n14591;
  assign n14593 = ~n7751 & ~n7869;
  assign n14594 = ~n8346 & n14593;
  assign n14595 = ~n9485 & n14594;
  assign n14596 = ~n10741 & n14595;
  assign n14597 = ~n12158 & n14596;
  assign n14598 = ~n13693 & n14597;
  assign n14599 = ~n9824 & ~n9929;
  assign n14600 = ~n11266 & n14599;
  assign n14601 = ~n11588 & n14600;
  assign n14602 = ~n13859 & n14601;
  assign n14603 = ~n14598 & ~n14602;
  assign n14604 = ~n14592 & n14603;
  assign n14605 = ~n3739 & ~n3940;
  assign n14606 = ~n4001 & n14605;
  assign n14607 = ~n5043 & n14606;
  assign n14608 = ~n5943 & n14607;
  assign n14609 = ~n6951 & n14608;
  assign n14610 = ~n8037 & n14609;
  assign n14611 = ~n9200 & n14610;
  assign n14612 = ~n10445 & n14611;
  assign n14613 = ~n11846 & n14612;
  assign n14614 = ~n13393 & n14613;
  assign n14615 = ~n2424 & ~n3066;
  assign n14616 = ~n3983 & n14615;
  assign n14617 = ~n4024 & n14616;
  assign n14618 = ~n4999 & n14617;
  assign n14619 = ~n5827 & n14618;
  assign n14620 = ~n6893 & n14619;
  assign n14621 = ~n7890 & n14620;
  assign n14622 = ~n9131 & n14621;
  assign n14623 = ~n10278 & n14622;
  assign n14624 = ~n11662 & n14623;
  assign n14625 = ~n13191 & n14624;
  assign n14626 = ~n14614 & ~n14625;
  assign n14627 = ~n6522 & ~n6784;
  assign n14628 = ~n7158 & n14627;
  assign n14629 = ~n8250 & n14628;
  assign n14630 = ~n9414 & n14629;
  assign n14631 = ~n10667 & n14630;
  assign n14632 = ~n12083 & n14631;
  assign n14633 = ~n13644 & n14632;
  assign n14634 = n3070 & n3072;
  assign n14635 = ~n2242 & n14634;
  assign n14636 = ~n3095 & n14635;
  assign n14637 = ~n3997 & n14636;
  assign n14638 = ~n4003 & n14637;
  assign n14639 = ~n4837 & n14638;
  assign n14640 = ~n5822 & n14639;
  assign n14641 = ~n6820 & n14640;
  assign n14642 = ~n7785 & n14641;
  assign n14643 = ~n9027 & n14642;
  assign n14644 = ~n10245 & n14643;
  assign n14645 = ~n13258 & n14644;
  assign n14646 = ~n13257 & n14645;
  assign n14647 = ~n11536 & n14646;
  assign n14648 = ~n13256 & n14647;
  assign n14649 = ~n13036 & n14648;
  assign n14650 = ~n13255 & n14649;
  assign n14651 = n13281 & n14650;
  assign n14652 = n13254 & n14651;
  assign n14653 = n13306 & n14652;
  assign n14654 = ~n1679 & ~n2242;
  assign n14655 = ~n3095 & n14654;
  assign n14656 = ~n3997 & n14655;
  assign n14657 = ~n4837 & n14656;
  assign n14658 = ~n5822 & n14657;
  assign n14659 = ~n6820 & n14658;
  assign n14660 = ~n7785 & n14659;
  assign n14661 = ~n9027 & n14660;
  assign n14662 = ~n10245 & n14661;
  assign n14663 = ~n11536 & n14662;
  assign n14664 = ~n13036 & n14663;
  assign n14665 = ~n14653 & n14664;
  assign n14666 = ~n14633 & ~n14665;
  assign n14667 = n14626 & n14666;
  assign n14668 = ~n8543 & ~n8834;
  assign n14669 = ~n10002 & n14668;
  assign n14670 = ~n11297 & n14669;
  assign n14671 = ~n12240 & n14670;
  assign n14672 = ~n13135 & n14671;
  assign n14673 = ~n12811 & ~n12902;
  assign n14674 = ~n14009 & n14673;
  assign n14675 = ~n14672 & ~n14674;
  assign n14676 = ~n12946 & ~n13093;
  assign n14677 = n719 & n781;
  assign n14678 = n1239 & n14677;
  assign n14679 = ~n1372 & n14678;
  assign n14680 = ~n2243 & n14679;
  assign n14681 = ~n3104 & n14680;
  assign n14682 = ~n3837 & n14681;
  assign n14683 = ~n3971 & n14682;
  assign n14684 = ~n4872 & n14683;
  assign n14685 = ~n5801 & n14684;
  assign n14686 = ~n6739 & n14685;
  assign n14687 = ~n7807 & n14686;
  assign n14688 = ~n8989 & n14687;
  assign n14689 = ~n10273 & n14688;
  assign n14690 = ~n13200 & n14689;
  assign n14691 = ~n13199 & n14690;
  assign n14692 = ~n11499 & n14691;
  assign n14693 = ~n13198 & n14692;
  assign n14694 = ~n13076 & n14693;
  assign n14695 = ~n13197 & n14694;
  assign n14696 = n13223 & n14695;
  assign n14697 = n13196 & n14696;
  assign n14698 = n13248 & n14697;
  assign n14699 = ~n688 & ~n1372;
  assign n14700 = ~n2243 & n14699;
  assign n14701 = ~n3104 & n14700;
  assign n14702 = ~n3971 & n14701;
  assign n14703 = ~n4872 & n14702;
  assign n14704 = ~n5801 & n14703;
  assign n14705 = ~n6739 & n14704;
  assign n14706 = ~n7807 & n14705;
  assign n14707 = ~n8989 & n14706;
  assign n14708 = ~n10273 & n14707;
  assign n14709 = ~n11499 & n14708;
  assign n14710 = ~n13076 & n14709;
  assign n14711 = ~n14698 & n14710;
  assign n14712 = ~n14676 & ~n14711;
  assign n14713 = n14675 & n14712;
  assign n14714 = n14667 & n14713;
  assign n14715 = n14604 & n14714;
  assign n14716 = n14583 & n14715;
  assign n14717 = ~n13393 & n13816;
  assign n14718 = ~n13135 & n13813;
  assign n14719 = ~n14717 & ~n14718;
  assign n14720 = ~n13558 & n13808;
  assign n14721 = ~n13644 & n13801;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = n14719 & n14722;
  assign n14724 = ~n13191 & n13815;
  assign n14725 = ~n13693 & n13805;
  assign n14726 = ~n14724 & ~n14725;
  assign n14727 = n13809 & ~n14698;
  assign n14728 = n13806 & ~n14653;
  assign n14729 = ~n14727 & ~n14728;
  assign n14730 = n14726 & n14729;
  assign n14731 = n13053 & ~n14467;
  assign n14732 = ~n13820 & n14731;
  assign n14733 = ~n14454 & n14732;
  assign n14734 = ~n14455 & n14733;
  assign n14735 = ~n13479 & n13812;
  assign n14736 = ~n14466 & ~n14572;
  assign n14737 = ~n14573 & n14736;
  assign n14738 = ~n14735 & n14737;
  assign n14739 = n14734 & n14738;
  assign n14740 = n14730 & n14739;
  assign n14741 = n14723 & n14740;
  assign n14742 = n13122 & ~n13820;
  assign n14743 = n13123 & ~n13906;
  assign n14744 = ~n14455 & ~n14743;
  assign n14745 = ~n14742 & n14744;
  assign n14746 = n8543 & ~n14568;
  assign n14747 = n8514 & ~n14519;
  assign n14748 = pi017 & ~n8574;
  assign n14749 = ~n8484 & n11377;
  assign n14750 = n14748 & n14749;
  assign n14751 = ~n8834 & n14750;
  assign n14752 = ~n10002 & n14751;
  assign n14753 = ~n14747 & n14752;
  assign n14754 = ~n14746 & n14753;
  assign n14755 = ~n11297 & n14754;
  assign n14756 = ~n12240 & n14755;
  assign n14757 = ~n14467 & n14756;
  assign n14758 = ~n14466 & n14757;
  assign n14759 = n14574 & n14758;
  assign n14760 = ~n13135 & ~n14454;
  assign n14761 = n14759 & n14760;
  assign n14762 = n13115 & ~n14073;
  assign n14763 = n13120 & ~n13479;
  assign n14764 = ~n14762 & ~n14763;
  assign n14765 = n14761 & n14764;
  assign n14766 = n14745 & n14765;
  assign n14767 = ~n13093 & n13096;
  assign n14768 = n13129 & ~n13393;
  assign n14769 = n13119 & ~n14698;
  assign n14770 = ~n14768 & ~n14769;
  assign n14771 = ~n14767 & n14770;
  assign n14772 = n13127 & ~n13693;
  assign n14773 = n13112 & ~n13644;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = n13116 & ~n14045;
  assign n14776 = n13126 & ~n13191;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = n14774 & n14777;
  assign n14779 = n13113 & ~n14653;
  assign n14780 = n13097 & ~n14009;
  assign n14781 = ~n14779 & ~n14780;
  assign n14782 = n13108 & ~n13859;
  assign n14783 = n13130 & ~n13558;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = n14781 & n14784;
  assign n14786 = n14778 & n14785;
  assign n14787 = n14771 & n14786;
  assign n14788 = n14766 & n14787;
  assign n14789 = n13183 & ~n13820;
  assign n14790 = n13169 & ~n13764;
  assign n14791 = n13172 & ~n13726;
  assign n14792 = ~n14790 & ~n14791;
  assign n14793 = ~n14789 & n14792;
  assign n14794 = n13136 & ~n13407;
  assign n14795 = n13142 & ~n13318;
  assign n14796 = n2631 & ~n14519;
  assign n14797 = n2424 & ~n14568;
  assign n14798 = ~n2602 & ~n2783;
  assign n14799 = n2573 & n14798;
  assign n14800 = ~n3066 & n14799;
  assign n14801 = ~n3983 & n14800;
  assign n14802 = ~n4003 & n14801;
  assign n14803 = ~n4024 & n14802;
  assign n14804 = ~n4999 & n14803;
  assign n14805 = ~n5827 & n14804;
  assign n14806 = ~n6893 & n14805;
  assign n14807 = ~n7890 & n14806;
  assign n14808 = ~n9131 & n14807;
  assign n14809 = ~n14797 & n14808;
  assign n14810 = ~n14796 & n14809;
  assign n14811 = ~n10278 & n14810;
  assign n14812 = ~n11662 & n14811;
  assign n14813 = ~n14795 & n14812;
  assign n14814 = ~n14794 & n14813;
  assign n14815 = n13138 & ~n13493;
  assign n14816 = n13137 & ~n13579;
  assign n14817 = ~n14815 & ~n14816;
  assign n14818 = n14814 & n14817;
  assign n14819 = n13171 & ~n13906;
  assign n14820 = ~n13191 & ~n14819;
  assign n14821 = n14818 & n14820;
  assign n14822 = n13186 & ~n14653;
  assign n14823 = n13144 & ~n14009;
  assign n14824 = ~n14822 & ~n14823;
  assign n14825 = n14821 & n14824;
  assign n14826 = n14793 & n14825;
  assign n14827 = ~n13093 & n13143;
  assign n14828 = n13179 & ~n13859;
  assign n14829 = n13164 & ~n14698;
  assign n14830 = ~n14828 & ~n14829;
  assign n14831 = ~n14827 & n14830;
  assign n14832 = n13176 & ~n14073;
  assign n14833 = n13168 & ~n13693;
  assign n14834 = ~n14832 & ~n14833;
  assign n14835 = n13141 & ~n14045;
  assign n14836 = n13185 & ~n13558;
  assign n14837 = ~n14835 & ~n14836;
  assign n14838 = n14834 & n14837;
  assign n14839 = ~n13135 & n13175;
  assign n14840 = n13182 & ~n13479;
  assign n14841 = ~n14839 & ~n14840;
  assign n14842 = n13163 & ~n13644;
  assign n14843 = n13178 & ~n13393;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = n14841 & n14844;
  assign n14846 = n14838 & n14845;
  assign n14847 = n14831 & n14846;
  assign n14848 = n14826 & n14847;
  assign n14849 = n13230 & ~n13726;
  assign n14850 = n13197 & ~n13820;
  assign n14851 = n13227 & ~n13764;
  assign n14852 = ~n14850 & ~n14851;
  assign n14853 = ~n14849 & n14852;
  assign n14854 = n13194 & ~n13493;
  assign n14855 = n13198 & ~n13318;
  assign n14856 = n688 & ~n14568;
  assign n14857 = n718 & ~n14519;
  assign n14858 = ~n780 & n4920;
  assign n14859 = n10294 & n14858;
  assign n14860 = ~n1372 & n14859;
  assign n14861 = ~n2243 & n14860;
  assign n14862 = ~n3104 & n14861;
  assign n14863 = ~n3971 & n14862;
  assign n14864 = ~n4003 & n14863;
  assign n14865 = ~n4872 & n14864;
  assign n14866 = ~n5801 & n14865;
  assign n14867 = ~n6739 & n14866;
  assign n14868 = ~n7807 & n14867;
  assign n14869 = ~n8989 & n14868;
  assign n14870 = ~n10273 & n14869;
  assign n14871 = ~n14857 & n14870;
  assign n14872 = ~n14856 & n14871;
  assign n14873 = ~n11499 & n14872;
  assign n14874 = ~n13076 & n14873;
  assign n14875 = ~n14855 & n14874;
  assign n14876 = ~n14854 & n14875;
  assign n14877 = n13193 & ~n13579;
  assign n14878 = n13192 & ~n13407;
  assign n14879 = ~n14877 & ~n14878;
  assign n14880 = n14876 & n14879;
  assign n14881 = n13229 & ~n13906;
  assign n14882 = ~n14698 & ~n14881;
  assign n14883 = n14880 & n14882;
  assign n14884 = n13240 & ~n14073;
  assign n14885 = n13243 & ~n13479;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = n14883 & n14886;
  assign n14888 = n14853 & n14887;
  assign n14889 = ~n13093 & n13200;
  assign n14890 = n13233 & ~n14653;
  assign n14891 = n13199 & ~n14009;
  assign n14892 = ~n14890 & ~n14891;
  assign n14893 = ~n14889 & n14892;
  assign n14894 = n13222 & ~n13393;
  assign n14895 = ~n13191 & n13236;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = n13241 & ~n14045;
  assign n14898 = n13244 & ~n13693;
  assign n14899 = ~n14897 & ~n14898;
  assign n14900 = n14896 & n14899;
  assign n14901 = n13226 & ~n13644;
  assign n14902 = n13234 & ~n13859;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n13135 & n13237;
  assign n14905 = n13221 & ~n13558;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = n14903 & n14906;
  assign n14908 = n14900 & n14907;
  assign n14909 = n14893 & n14908;
  assign n14910 = n14888 & n14909;
  assign n14911 = n13288 & ~n13726;
  assign n14912 = n13287 & ~n13906;
  assign n14913 = n13285 & ~n13764;
  assign n14914 = ~n14912 & ~n14913;
  assign n14915 = ~n14911 & n14914;
  assign n14916 = n13251 & ~n13579;
  assign n14917 = n13256 & ~n13318;
  assign n14918 = n1679 & ~n14568;
  assign n14919 = n1710 & ~n14519;
  assign n14920 = pi003 & ~n1740;
  assign n14921 = n13259 & n14920;
  assign n14922 = ~n2242 & n14921;
  assign n14923 = ~n3095 & n14922;
  assign n14924 = ~n3997 & n14923;
  assign n14925 = ~n4003 & n14924;
  assign n14926 = ~n4837 & n14925;
  assign n14927 = ~n5822 & n14926;
  assign n14928 = ~n6820 & n14927;
  assign n14929 = ~n7785 & n14928;
  assign n14930 = ~n9027 & n14929;
  assign n14931 = ~n10245 & n14930;
  assign n14932 = ~n14919 & n14931;
  assign n14933 = ~n14918 & n14932;
  assign n14934 = ~n11536 & n14933;
  assign n14935 = ~n13036 & n14934;
  assign n14936 = ~n14917 & n14935;
  assign n14937 = ~n14916 & n14936;
  assign n14938 = n13250 & ~n13407;
  assign n14939 = n13252 & ~n13493;
  assign n14940 = ~n14938 & ~n14939;
  assign n14941 = n14937 & n14940;
  assign n14942 = n13294 & ~n13820;
  assign n14943 = ~n14653 & ~n14942;
  assign n14944 = n14941 & n14943;
  assign n14945 = n13295 & ~n13859;
  assign n14946 = n13301 & ~n13644;
  assign n14947 = ~n14945 & ~n14946;
  assign n14948 = n14944 & n14947;
  assign n14949 = n14915 & n14948;
  assign n14950 = ~n13093 & n13258;
  assign n14951 = n13302 & ~n13693;
  assign n14952 = n13298 & ~n14698;
  assign n14953 = ~n14951 & ~n14952;
  assign n14954 = ~n14950 & n14953;
  assign n14955 = ~n13135 & n13299;
  assign n14956 = n13292 & ~n13393;
  assign n14957 = ~n14955 & ~n14956;
  assign n14958 = n13279 & ~n14045;
  assign n14959 = n13280 & ~n13558;
  assign n14960 = ~n14958 & ~n14959;
  assign n14961 = n14957 & n14960;
  assign n14962 = n13257 & ~n14009;
  assign n14963 = n13255 & ~n14073;
  assign n14964 = ~n14962 & ~n14963;
  assign n14965 = n13291 & ~n13479;
  assign n14966 = ~n13191 & n13284;
  assign n14967 = ~n14965 & ~n14966;
  assign n14968 = n14964 & n14967;
  assign n14969 = n14961 & n14968;
  assign n14970 = n14954 & n14969;
  assign n14971 = n14949 & n14970;
  assign n14972 = ~n14910 & ~n14971;
  assign n14973 = ~n14848 & n14972;
  assign n14974 = n13316 & ~n14698;
  assign n14975 = n13313 & ~n13318;
  assign n14976 = ~n14974 & n14975;
  assign n14977 = ~n13191 & n13315;
  assign n14978 = n13310 & ~n14653;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = n14976 & n14979;
  assign n14981 = ~n2783 & n3846;
  assign n14982 = n7972 & n14981;
  assign n14983 = ~n3066 & n14982;
  assign n14984 = ~n3983 & n14983;
  assign n14985 = ~n4003 & n14984;
  assign n14986 = ~n4024 & n14985;
  assign n14987 = ~n4999 & n14986;
  assign n14988 = ~n5827 & n14987;
  assign n14989 = ~n6893 & n14988;
  assign n14990 = ~n7890 & n14989;
  assign n14991 = ~n9131 & n14990;
  assign n14992 = ~n14797 & n14991;
  assign n14993 = ~n14796 & n14992;
  assign n14994 = ~n10278 & n14993;
  assign n14995 = ~n11662 & n14994;
  assign n14996 = ~n14795 & n14995;
  assign n14997 = ~n14794 & n14996;
  assign n14998 = n14817 & n14997;
  assign n14999 = n14820 & n14998;
  assign n15000 = n14824 & n14999;
  assign n15001 = n14793 & n15000;
  assign n15002 = n14847 & n15001;
  assign n15003 = ~n14980 & ~n15002;
  assign n15004 = ~n14973 & n15003;
  assign n15005 = n13373 & ~n13726;
  assign n15006 = n13374 & ~n13764;
  assign n15007 = n13384 & ~n13820;
  assign n15008 = ~n15006 & ~n15007;
  assign n15009 = ~n15005 & n15008;
  assign n15010 = n13342 & ~n13407;
  assign n15011 = n3739 & ~n14568;
  assign n15012 = n3769 & ~n14519;
  assign n15013 = ~n3591 & ~n3710;
  assign n15014 = n4103 & n15013;
  assign n15015 = ~n3940 & n15014;
  assign n15016 = ~n4001 & n15015;
  assign n15017 = ~n5043 & n15016;
  assign n15018 = ~n5943 & n15017;
  assign n15019 = ~n6951 & n15018;
  assign n15020 = ~n8037 & n15019;
  assign n15021 = ~n9200 & n15020;
  assign n15022 = ~n15012 & n15021;
  assign n15023 = ~n15011 & n15022;
  assign n15024 = ~n10445 & n15023;
  assign n15025 = ~n11846 & n15024;
  assign n15026 = ~n14467 & n15025;
  assign n15027 = ~n15010 & n15026;
  assign n15028 = n13341 & ~n13493;
  assign n15029 = n13343 & ~n13579;
  assign n15030 = ~n15028 & ~n15029;
  assign n15031 = n15027 & n15030;
  assign n15032 = n13377 & ~n13906;
  assign n15033 = ~n13393 & ~n15032;
  assign n15034 = n15031 & n15033;
  assign n15035 = n13370 & ~n13479;
  assign n15036 = n13378 & ~n13693;
  assign n15037 = ~n15035 & ~n15036;
  assign n15038 = n15034 & n15037;
  assign n15039 = n15009 & n15038;
  assign n15040 = ~n13093 & n13348;
  assign n15041 = ~n13191 & n13380;
  assign n15042 = n13365 & ~n14698;
  assign n15043 = ~n15041 & ~n15042;
  assign n15044 = ~n15040 & n15043;
  assign n15045 = n13387 & ~n14653;
  assign n15046 = n13366 & ~n13558;
  assign n15047 = ~n15045 & ~n15046;
  assign n15048 = n13371 & ~n14045;
  assign n15049 = n13346 & ~n13644;
  assign n15050 = ~n15048 & ~n15049;
  assign n15051 = n15047 & n15050;
  assign n15052 = ~n13135 & n13388;
  assign n15053 = n13385 & ~n14073;
  assign n15054 = ~n15052 & ~n15053;
  assign n15055 = n13381 & ~n13859;
  assign n15056 = n13347 & ~n14009;
  assign n15057 = ~n15055 & ~n15056;
  assign n15058 = n15054 & n15057;
  assign n15059 = n15051 & n15058;
  assign n15060 = n15044 & n15059;
  assign n15061 = n15039 & n15060;
  assign n15062 = ~n13318 & n13394;
  assign n15063 = ~n14974 & n15062;
  assign n15064 = n14979 & n15063;
  assign n15065 = ~n15061 & ~n15064;
  assign n15066 = ~n15004 & n15065;
  assign n15067 = n13404 & ~n14653;
  assign n15068 = ~n14467 & n14573;
  assign n15069 = ~n15067 & n15068;
  assign n15070 = n13403 & ~n14698;
  assign n15071 = ~n13393 & n13402;
  assign n15072 = ~n13191 & n13399;
  assign n15073 = ~n15071 & ~n15072;
  assign n15074 = ~n15070 & n15073;
  assign n15075 = n15069 & n15074;
  assign n15076 = n10461 & n13408;
  assign n15077 = ~n3940 & n15076;
  assign n15078 = ~n4001 & n15077;
  assign n15079 = ~n5043 & n15078;
  assign n15080 = ~n5943 & n15079;
  assign n15081 = ~n6951 & n15080;
  assign n15082 = ~n8037 & n15081;
  assign n15083 = ~n9200 & n15082;
  assign n15084 = ~n15012 & n15083;
  assign n15085 = ~n15011 & n15084;
  assign n15086 = ~n10445 & n15085;
  assign n15087 = ~n11846 & n15086;
  assign n15088 = ~n14467 & n15087;
  assign n15089 = ~n15010 & n15088;
  assign n15090 = n15030 & n15089;
  assign n15091 = n15033 & n15090;
  assign n15092 = n15037 & n15091;
  assign n15093 = n15009 & n15092;
  assign n15094 = n15060 & n15093;
  assign n15095 = ~n15075 & ~n15094;
  assign n15096 = ~n15066 & n15095;
  assign n15097 = ~n13407 & n13428;
  assign n15098 = ~n14467 & n15097;
  assign n15099 = ~n15067 & n15098;
  assign n15100 = n15074 & n15099;
  assign n15101 = n13457 & ~n13764;
  assign n15102 = n13471 & ~n13820;
  assign n15103 = n13460 & ~n13726;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = ~n15101 & n15104;
  assign n15106 = n4736 & ~n14519;
  assign n15107 = n4707 & ~n14568;
  assign n15108 = n4491 & ~n4817;
  assign n15109 = ~n4902 & n15108;
  assign n15110 = ~n6001 & n15109;
  assign n15111 = ~n7014 & n15110;
  assign n15112 = ~n8114 & n15111;
  assign n15113 = ~n9276 & n15112;
  assign n15114 = ~n15107 & n15113;
  assign n15115 = ~n15106 & n15114;
  assign n15116 = ~n10523 & n15115;
  assign n15117 = ~n11928 & n15116;
  assign n15118 = ~n14467 & n15117;
  assign n15119 = ~n14573 & n15118;
  assign n15120 = n13433 & ~n13493;
  assign n15121 = n13432 & ~n13579;
  assign n15122 = ~n15120 & ~n15121;
  assign n15123 = n15119 & n15122;
  assign n15124 = n13459 & ~n13906;
  assign n15125 = ~n13479 & ~n15124;
  assign n15126 = n15123 & n15125;
  assign n15127 = n13463 & ~n14073;
  assign n15128 = n13456 & ~n13693;
  assign n15129 = ~n15127 & ~n15128;
  assign n15130 = n15126 & n15129;
  assign n15131 = n15105 & n15130;
  assign n15132 = ~n13093 & n13438;
  assign n15133 = n13470 & ~n13558;
  assign n15134 = n13452 & ~n14698;
  assign n15135 = ~n15133 & ~n15134;
  assign n15136 = ~n15132 & n15135;
  assign n15137 = n13464 & ~n13859;
  assign n15138 = ~n13393 & n13466;
  assign n15139 = ~n15137 & ~n15138;
  assign n15140 = n13436 & ~n14045;
  assign n15141 = ~n13191 & n13451;
  assign n15142 = ~n15140 & ~n15141;
  assign n15143 = n15139 & n15142;
  assign n15144 = n13474 & ~n14653;
  assign n15145 = n13437 & ~n14009;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = n13467 & ~n13644;
  assign n15148 = ~n13135 & n13473;
  assign n15149 = ~n15147 & ~n15148;
  assign n15150 = n15146 & n15149;
  assign n15151 = n15143 & n15150;
  assign n15152 = n15136 & n15151;
  assign n15153 = n15131 & n15152;
  assign n15154 = ~n15100 & ~n15153;
  assign n15155 = ~n15096 & n15154;
  assign n15156 = n13489 & ~n14653;
  assign n15157 = ~n14467 & n14572;
  assign n15158 = ~n14573 & n15157;
  assign n15159 = ~n15156 & n15158;
  assign n15160 = n13484 & ~n14698;
  assign n15161 = ~n13479 & n13482;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = ~n13393 & n13490;
  assign n15164 = ~n13191 & n13483;
  assign n15165 = ~n15163 & ~n15164;
  assign n15166 = n15162 & n15165;
  assign n15167 = n15159 & n15166;
  assign n15168 = ~pi009 & ~n4401;
  assign n15169 = n13494 & n15168;
  assign n15170 = ~n4817 & n15169;
  assign n15171 = ~n4902 & n15170;
  assign n15172 = ~n6001 & n15171;
  assign n15173 = ~n7014 & n15172;
  assign n15174 = ~n8114 & n15173;
  assign n15175 = ~n9276 & n15174;
  assign n15176 = ~n15107 & n15175;
  assign n15177 = ~n15106 & n15176;
  assign n15178 = ~n10523 & n15177;
  assign n15179 = ~n11928 & n15178;
  assign n15180 = ~n14467 & n15179;
  assign n15181 = ~n14573 & n15180;
  assign n15182 = n15122 & n15181;
  assign n15183 = n15125 & n15182;
  assign n15184 = n15129 & n15183;
  assign n15185 = n15105 & n15184;
  assign n15186 = n15152 & n15185;
  assign n15187 = ~n15167 & ~n15186;
  assign n15188 = ~n15155 & n15187;
  assign n15189 = n13550 & ~n13820;
  assign n15190 = n13536 & ~n13764;
  assign n15191 = n13539 & ~n13726;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = ~n15189 & n15192;
  assign n15194 = n5408 & ~n14519;
  assign n15195 = n5378 & ~n14568;
  assign n15196 = ~n5808 & n7096;
  assign n15197 = ~n6056 & n15196;
  assign n15198 = ~n7073 & n15197;
  assign n15199 = ~n8179 & n15198;
  assign n15200 = ~n9344 & n15199;
  assign n15201 = ~n15195 & n15200;
  assign n15202 = ~n15194 & n15201;
  assign n15203 = ~n10594 & n15202;
  assign n15204 = ~n12005 & n15203;
  assign n15205 = ~n14467 & n15204;
  assign n15206 = ~n14572 & n15205;
  assign n15207 = n13513 & ~n13579;
  assign n15208 = ~n14573 & ~n15207;
  assign n15209 = n15206 & n15208;
  assign n15210 = n13538 & ~n13906;
  assign n15211 = ~n13558 & ~n15210;
  assign n15212 = n15209 & n15211;
  assign n15213 = n13543 & ~n13859;
  assign n15214 = n13553 & ~n14653;
  assign n15215 = ~n15213 & ~n15214;
  assign n15216 = n15212 & n15215;
  assign n15217 = n15193 & n15216;
  assign n15218 = ~n13093 & n13517;
  assign n15219 = ~n13393 & n13545;
  assign n15220 = n13531 & ~n14698;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = ~n15218 & n15221;
  assign n15223 = n13542 & ~n14073;
  assign n15224 = n13535 & ~n13693;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = n13515 & ~n14045;
  assign n15227 = n13546 & ~n13644;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = n15225 & n15228;
  assign n15230 = ~n13135 & n13552;
  assign n15231 = n13516 & ~n14009;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = ~n13191 & n13530;
  assign n15234 = ~n13479 & n13549;
  assign n15235 = ~n15233 & ~n15234;
  assign n15236 = n15232 & n15235;
  assign n15237 = n15229 & n15236;
  assign n15238 = n15222 & n15237;
  assign n15239 = n15217 & n15238;
  assign n15240 = ~n13493 & n13559;
  assign n15241 = ~n14467 & n15240;
  assign n15242 = ~n14573 & n15241;
  assign n15243 = ~n15156 & n15242;
  assign n15244 = n15166 & n15243;
  assign n15245 = ~n15239 & ~n15244;
  assign n15246 = ~n15188 & n15245;
  assign n15247 = ~n5349 & n5687;
  assign n15248 = n13581 & n15247;
  assign n15249 = ~n5808 & n15248;
  assign n15250 = ~n6056 & n15249;
  assign n15251 = ~n7073 & n15250;
  assign n15252 = ~n8179 & n15251;
  assign n15253 = ~n9344 & n15252;
  assign n15254 = ~n15195 & n15253;
  assign n15255 = ~n15194 & n15254;
  assign n15256 = ~n10594 & n15255;
  assign n15257 = ~n12005 & n15256;
  assign n15258 = ~n14467 & n15257;
  assign n15259 = ~n14572 & n15258;
  assign n15260 = n15208 & n15259;
  assign n15261 = n15211 & n15260;
  assign n15262 = n15215 & n15261;
  assign n15263 = n15193 & n15262;
  assign n15264 = n15238 & n15263;
  assign n15265 = ~n13191 & n13570;
  assign n15266 = n13576 & ~n14653;
  assign n15267 = n13575 & ~n14698;
  assign n15268 = ~n15266 & ~n15267;
  assign n15269 = ~n15265 & n15268;
  assign n15270 = ~n13479 & n13569;
  assign n15271 = n14466 & ~n14467;
  assign n15272 = n14574 & n15271;
  assign n15273 = ~n15270 & n15272;
  assign n15274 = ~n13393 & n13567;
  assign n15275 = ~n13558 & n13566;
  assign n15276 = ~n15274 & ~n15275;
  assign n15277 = n15273 & n15276;
  assign n15278 = n15269 & n15277;
  assign n15279 = ~n15264 & ~n15278;
  assign n15280 = ~n15246 & n15279;
  assign n15281 = n13622 & ~n13726;
  assign n15282 = n13625 & ~n13764;
  assign n15283 = n13635 & ~n13820;
  assign n15284 = ~n15282 & ~n15283;
  assign n15285 = ~n15281 & n15284;
  assign n15286 = n6522 & ~n14568;
  assign n15287 = n6613 & ~n14519;
  assign n15288 = ~n6584 & ~n6643;
  assign n15289 = n12054 & n15288;
  assign n15290 = ~n6784 & n15289;
  assign n15291 = ~n7158 & n15290;
  assign n15292 = ~n8250 & n15291;
  assign n15293 = ~n9414 & n15292;
  assign n15294 = ~n15287 & n15293;
  assign n15295 = ~n15286 & n15294;
  assign n15296 = ~n10667 & n15295;
  assign n15297 = ~n12083 & n15296;
  assign n15298 = ~n14467 & n15297;
  assign n15299 = ~n14466 & n15298;
  assign n15300 = n14574 & n15299;
  assign n15301 = n13628 & ~n13906;
  assign n15302 = ~n13644 & ~n15301;
  assign n15303 = n15300 & n15302;
  assign n15304 = n13601 & ~n14009;
  assign n15305 = n13638 & ~n14653;
  assign n15306 = ~n15304 & ~n15305;
  assign n15307 = n15303 & n15306;
  assign n15308 = n15285 & n15307;
  assign n15309 = ~n13093 & n13602;
  assign n15310 = n13629 & ~n13859;
  assign n15311 = n13616 & ~n14698;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = ~n15309 & n15312;
  assign n15314 = n13636 & ~n14073;
  assign n15315 = ~n13558 & n13600;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = n13624 & ~n14045;
  assign n15318 = n13621 & ~n13693;
  assign n15319 = ~n15317 & ~n15318;
  assign n15320 = n15316 & n15319;
  assign n15321 = ~n13191 & n13631;
  assign n15322 = ~n13479 & n13639;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n13135 & n13632;
  assign n15325 = ~n13393 & n13617;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = n15323 & n15326;
  assign n15328 = n15320 & n15327;
  assign n15329 = n15313 & n15328;
  assign n15330 = n15308 & n15329;
  assign n15331 = ~n13579 & n13645;
  assign n15332 = ~n14467 & n15331;
  assign n15333 = n14574 & n15332;
  assign n15334 = ~n15270 & n15333;
  assign n15335 = n15276 & n15334;
  assign n15336 = n15269 & n15335;
  assign n15337 = ~n15330 & ~n15336;
  assign n15338 = ~n15280 & n15337;
  assign n15339 = n13673 & ~n13764;
  assign n15340 = n13674 & ~n13906;
  assign n15341 = n13678 & ~n13820;
  assign n15342 = ~n15340 & ~n15341;
  assign n15343 = ~n15339 & n15342;
  assign n15344 = n7751 & ~n14568;
  assign n15345 = n7722 & ~n14519;
  assign n15346 = n7693 & n8364;
  assign n15347 = ~n7869 & n15346;
  assign n15348 = ~n8346 & n15347;
  assign n15349 = ~n9485 & n15348;
  assign n15350 = ~n15345 & n15349;
  assign n15351 = ~n15344 & n15350;
  assign n15352 = ~n10741 & n15351;
  assign n15353 = ~n12158 & n15352;
  assign n15354 = ~n14467 & n15353;
  assign n15355 = ~n14466 & n15354;
  assign n15356 = n14574 & n15355;
  assign n15357 = ~n13693 & ~n14455;
  assign n15358 = n15356 & n15357;
  assign n15359 = n13665 & ~n14073;
  assign n15360 = ~n13479 & n13677;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = n15358 & n15361;
  assign n15363 = n15343 & n15362;
  assign n15364 = ~n13093 & n13652;
  assign n15365 = ~n13393 & n13685;
  assign n15366 = n13688 & ~n14698;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~n15364 & n15367;
  assign n15369 = ~n13644 & n13681;
  assign n15370 = ~n13135 & n13684;
  assign n15371 = ~n15369 & ~n15370;
  assign n15372 = n13680 & ~n14045;
  assign n15373 = ~n13191 & n13666;
  assign n15374 = ~n15372 & ~n15373;
  assign n15375 = n15371 & n15374;
  assign n15376 = n13671 & ~n14653;
  assign n15377 = n13653 & ~n14009;
  assign n15378 = ~n15376 & ~n15377;
  assign n15379 = n13670 & ~n13859;
  assign n15380 = ~n13558 & n13687;
  assign n15381 = ~n15379 & ~n15380;
  assign n15382 = n15378 & n15381;
  assign n15383 = n15375 & n15382;
  assign n15384 = n15368 & n15383;
  assign n15385 = n15363 & n15384;
  assign n15386 = ~n6643 & n7175;
  assign n15387 = n10675 & n15386;
  assign n15388 = ~n6784 & n15387;
  assign n15389 = ~n7158 & n15388;
  assign n15390 = ~n8250 & n15389;
  assign n15391 = ~n9414 & n15390;
  assign n15392 = ~n15287 & n15391;
  assign n15393 = ~n15286 & n15392;
  assign n15394 = ~n10667 & n15393;
  assign n15395 = ~n12083 & n15394;
  assign n15396 = ~n14467 & n15395;
  assign n15397 = ~n14466 & n15396;
  assign n15398 = n14574 & n15397;
  assign n15399 = n15302 & n15398;
  assign n15400 = n15306 & n15399;
  assign n15401 = n15285 & n15400;
  assign n15402 = n15329 & n15401;
  assign n15403 = ~n13393 & n13721;
  assign n15404 = ~n13558 & n13722;
  assign n15405 = ~n13479 & n13711;
  assign n15406 = ~n15404 & ~n15405;
  assign n15407 = ~n15403 & n15406;
  assign n15408 = n13052 & ~n14467;
  assign n15409 = ~n13726 & n15408;
  assign n15410 = n14737 & n15409;
  assign n15411 = n13710 & ~n14698;
  assign n15412 = ~n13191 & n13713;
  assign n15413 = ~n15411 & ~n15412;
  assign n15414 = ~n13644 & n13714;
  assign n15415 = n13717 & ~n14653;
  assign n15416 = ~n15414 & ~n15415;
  assign n15417 = n15413 & n15416;
  assign n15418 = n15410 & n15417;
  assign n15419 = n15407 & n15418;
  assign n15420 = ~n15402 & ~n15419;
  assign n15421 = ~n15385 & n15420;
  assign n15422 = ~n15338 & n15421;
  assign n15423 = ~n7475 & ~n7692;
  assign n15424 = ~n7505 & n15423;
  assign n15425 = n8357 & n15424;
  assign n15426 = ~n7869 & n15425;
  assign n15427 = ~n8346 & n15426;
  assign n15428 = ~n9485 & n15427;
  assign n15429 = ~n15345 & n15428;
  assign n15430 = ~n15344 & n15429;
  assign n15431 = ~n10741 & n15430;
  assign n15432 = ~n12158 & n15431;
  assign n15433 = ~n14467 & n15432;
  assign n15434 = ~n14466 & n15433;
  assign n15435 = n14574 & n15434;
  assign n15436 = n15357 & n15435;
  assign n15437 = n15361 & n15436;
  assign n15438 = n15343 & n15437;
  assign n15439 = n15384 & n15438;
  assign n15440 = ~n12121 & n13765;
  assign n15441 = ~n14467 & n15440;
  assign n15442 = ~n13726 & n15441;
  assign n15443 = n14737 & n15442;
  assign n15444 = n15417 & n15443;
  assign n15445 = n15407 & n15444;
  assign n15446 = ~n13693 & n13749;
  assign n15447 = n13756 & ~n14698;
  assign n15448 = ~n15446 & ~n15447;
  assign n15449 = ~n13644 & n13748;
  assign n15450 = ~n13393 & n13753;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = n15448 & n15451;
  assign n15453 = n12973 & ~n14467;
  assign n15454 = ~n13764 & n15453;
  assign n15455 = ~n14455 & n15454;
  assign n15456 = n14737 & n15455;
  assign n15457 = ~n13191 & n13745;
  assign n15458 = ~n13479 & n13752;
  assign n15459 = ~n15457 & ~n15458;
  assign n15460 = ~n13558 & n13755;
  assign n15461 = n13746 & ~n14653;
  assign n15462 = ~n15460 & ~n15461;
  assign n15463 = n15459 & n15462;
  assign n15464 = n15456 & n15463;
  assign n15465 = n15452 & n15464;
  assign n15466 = ~n15445 & ~n15465;
  assign n15467 = ~n15439 & n15466;
  assign n15468 = ~n15422 & n15467;
  assign n15469 = n8485 & n13098;
  assign n15470 = ~n8834 & n15469;
  assign n15471 = ~n10002 & n15470;
  assign n15472 = ~n14747 & n15471;
  assign n15473 = ~n14746 & n15472;
  assign n15474 = ~n11297 & n15473;
  assign n15475 = ~n12240 & n15474;
  assign n15476 = ~n14467 & n15475;
  assign n15477 = ~n14466 & n15476;
  assign n15478 = n14574 & n15477;
  assign n15479 = n14760 & n15478;
  assign n15480 = n14764 & n15479;
  assign n15481 = n14745 & n15480;
  assign n15482 = n14787 & n15481;
  assign n15483 = ~n12181 & n13775;
  assign n15484 = ~n14467 & n15483;
  assign n15485 = ~n13764 & n15484;
  assign n15486 = ~n14455 & n15485;
  assign n15487 = n14737 & n15486;
  assign n15488 = n15463 & n15487;
  assign n15489 = n15452 & n15488;
  assign n15490 = ~n15482 & ~n15489;
  assign n15491 = ~n15468 & n15490;
  assign n15492 = ~n14788 & ~n15491;
  assign n15493 = ~n14741 & ~n15492;
  assign n15494 = n13851 & ~n13906;
  assign n15495 = n14456 & ~n15494;
  assign n15496 = n9824 & ~n14568;
  assign n15497 = n9717 & ~n14519;
  assign n15498 = ~n9793 & ~n9854;
  assign n15499 = n11562 & n15498;
  assign n15500 = ~n9929 & n15499;
  assign n15501 = ~n15497 & n15500;
  assign n15502 = ~n15496 & n15501;
  assign n15503 = ~n11266 & n15502;
  assign n15504 = ~n11588 & n15503;
  assign n15505 = ~n14467 & n15504;
  assign n15506 = ~n14466 & n15505;
  assign n15507 = n14574 & n15506;
  assign n15508 = ~n13859 & ~n14452;
  assign n15509 = n15507 & n15508;
  assign n15510 = n13824 & ~n14009;
  assign n15511 = ~n13693 & n13840;
  assign n15512 = ~n15510 & ~n15511;
  assign n15513 = n15509 & n15512;
  assign n15514 = n15495 & n15513;
  assign n15515 = ~n13093 & n13823;
  assign n15516 = ~n13558 & n13843;
  assign n15517 = n13844 & ~n14698;
  assign n15518 = ~n15516 & ~n15517;
  assign n15519 = ~n15515 & n15518;
  assign n15520 = ~n13135 & n13837;
  assign n15521 = ~n13191 & n13839;
  assign n15522 = ~n15520 & ~n15521;
  assign n15523 = ~n13479 & n13846;
  assign n15524 = n13850 & ~n14045;
  assign n15525 = ~n15523 & ~n15524;
  assign n15526 = n15522 & n15525;
  assign n15527 = n13853 & ~n14653;
  assign n15528 = ~n13644 & n13836;
  assign n15529 = ~n15527 & ~n15528;
  assign n15530 = ~n13393 & n13847;
  assign n15531 = n13854 & ~n14073;
  assign n15532 = ~n15530 & ~n15531;
  assign n15533 = n15529 & n15532;
  assign n15534 = n15526 & n15533;
  assign n15535 = n15519 & n15534;
  assign n15536 = n15514 & n15535;
  assign n15537 = ~n11611 & n13860;
  assign n15538 = ~n14467 & n15537;
  assign n15539 = ~n13820 & n15538;
  assign n15540 = ~n14454 & n15539;
  assign n15541 = ~n14455 & n15540;
  assign n15542 = n14738 & n15541;
  assign n15543 = n14730 & n15542;
  assign n15544 = n14723 & n15543;
  assign n15545 = ~n15536 & ~n15544;
  assign n15546 = ~n15493 & n15545;
  assign n15547 = ~pi019 & ~n9913;
  assign n15548 = n9794 & ~n9854;
  assign n15549 = n15547 & n15548;
  assign n15550 = ~n9929 & n15549;
  assign n15551 = ~n15497 & n15550;
  assign n15552 = ~n15496 & n15551;
  assign n15553 = ~n11266 & n15552;
  assign n15554 = ~n11588 & n15553;
  assign n15555 = ~n14467 & n15554;
  assign n15556 = ~n14466 & n15555;
  assign n15557 = n14574 & n15556;
  assign n15558 = n15508 & n15557;
  assign n15559 = n15512 & n15558;
  assign n15560 = n15495 & n15559;
  assign n15561 = n15535 & n15560;
  assign n15562 = n12972 & ~n14467;
  assign n15563 = ~n13906 & n15562;
  assign n15564 = ~n14452 & n15563;
  assign n15565 = n14456 & n15564;
  assign n15566 = ~n13479 & n13895;
  assign n15567 = n14737 & ~n15566;
  assign n15568 = ~n13693 & n13891;
  assign n15569 = ~n13644 & n13899;
  assign n15570 = ~n15568 & ~n15569;
  assign n15571 = n15567 & n15570;
  assign n15572 = n15565 & n15571;
  assign n15573 = ~n13191 & n13898;
  assign n15574 = n13883 & ~n14653;
  assign n15575 = ~n13135 & n13892;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = ~n15573 & n15576;
  assign n15578 = ~n13859 & n13882;
  assign n15579 = ~n13558 & n13901;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = n13894 & ~n14698;
  assign n15582 = ~n13393 & n13902;
  assign n15583 = ~n15581 & ~n15582;
  assign n15584 = n15580 & n15583;
  assign n15585 = n15577 & n15584;
  assign n15586 = n15572 & n15585;
  assign n15587 = ~n13693 & n14058;
  assign n15588 = ~n13393 & n14054;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = ~n13644 & n14051;
  assign n15591 = ~n13479 & n14068;
  assign n15592 = ~n15590 & ~n15591;
  assign n15593 = n15589 & n15592;
  assign n15594 = ~n14452 & ~n14454;
  assign n15595 = ~n14455 & n15594;
  assign n15596 = n13055 & ~n14467;
  assign n15597 = ~n14466 & n15596;
  assign n15598 = n14574 & n15597;
  assign n15599 = ~n14073 & ~n14451;
  assign n15600 = n15598 & n15599;
  assign n15601 = n15595 & n15600;
  assign n15602 = n15593 & n15601;
  assign n15603 = n14061 & ~n14653;
  assign n15604 = ~n13859 & n14062;
  assign n15605 = n14052 & ~n14698;
  assign n15606 = ~n15604 & ~n15605;
  assign n15607 = ~n15603 & n15606;
  assign n15608 = ~n13191 & n14065;
  assign n15609 = ~n13558 & n14059;
  assign n15610 = ~n15608 & ~n15609;
  assign n15611 = ~n13135 & n14067;
  assign n15612 = ~n14045 & n14055;
  assign n15613 = ~n15611 & ~n15612;
  assign n15614 = n15610 & n15613;
  assign n15615 = n15607 & n15614;
  assign n15616 = n15602 & n15615;
  assign n15617 = ~n15586 & ~n15616;
  assign n15618 = ~n15561 & n15617;
  assign n15619 = n11133 & ~n14568;
  assign n15620 = n10909 & ~n14519;
  assign n15621 = n12315 & n12317;
  assign n15622 = ~n11188 & n15621;
  assign n15623 = ~n15620 & n15622;
  assign n15624 = ~n15619 & n15623;
  assign n15625 = ~n12380 & n15624;
  assign n15626 = ~n14467 & n15625;
  assign n15627 = ~n14466 & n15626;
  assign n15628 = n14574 & n15627;
  assign n15629 = ~n14045 & ~n14451;
  assign n15630 = n15628 & n15629;
  assign n15631 = ~n13393 & n14026;
  assign n15632 = n14033 & ~n14653;
  assign n15633 = ~n15631 & ~n15632;
  assign n15634 = n15630 & n15633;
  assign n15635 = n15595 & n15634;
  assign n15636 = ~n13135 & n14023;
  assign n15637 = ~n13191 & n14040;
  assign n15638 = ~n13693 & n14030;
  assign n15639 = ~n15637 & ~n15638;
  assign n15640 = ~n15636 & n15639;
  assign n15641 = n14034 & ~n14698;
  assign n15642 = ~n13479 & n14024;
  assign n15643 = ~n15641 & ~n15642;
  assign n15644 = ~n14009 & n14011;
  assign n15645 = ~n13558 & n14027;
  assign n15646 = ~n15644 & ~n15645;
  assign n15647 = n15643 & n15646;
  assign n15648 = ~n13859 & n14039;
  assign n15649 = n14037 & ~n14073;
  assign n15650 = ~n15648 & ~n15649;
  assign n15651 = ~n13093 & n14010;
  assign n15652 = ~n13644 & n14031;
  assign n15653 = ~n15651 & ~n15652;
  assign n15654 = n15650 & n15653;
  assign n15655 = n15647 & n15654;
  assign n15656 = n15640 & n15655;
  assign n15657 = n15635 & n15656;
  assign n15658 = n12671 & ~n14519;
  assign n15659 = n12811 & ~n14568;
  assign n15660 = ~n12902 & n13912;
  assign n15661 = ~n15659 & n15660;
  assign n15662 = ~n15658 & n15661;
  assign n15663 = ~n14467 & n15662;
  assign n15664 = ~n14466 & n15663;
  assign n15665 = n14574 & n15664;
  assign n15666 = ~n14009 & ~n14451;
  assign n15667 = n15665 & n15666;
  assign n15668 = ~n13558 & n13949;
  assign n15669 = ~n14577 & ~n15668;
  assign n15670 = n15667 & n15669;
  assign n15671 = n15595 & n15670;
  assign n15672 = ~n13644 & n13990;
  assign n15673 = ~n13135 & n13982;
  assign n15674 = ~n13093 & n13908;
  assign n15675 = ~n15673 & ~n15674;
  assign n15676 = ~n15672 & n15675;
  assign n15677 = ~n13693 & n13978;
  assign n15678 = ~n13859 & n13933;
  assign n15679 = ~n15677 & ~n15678;
  assign n15680 = n13963 & ~n14698;
  assign n15681 = ~n13191 & n13930;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = n15679 & n15682;
  assign n15684 = ~n13479 & n13942;
  assign n15685 = ~n13393 & n13972;
  assign n15686 = ~n15684 & ~n15685;
  assign n15687 = n14004 & ~n14045;
  assign n15688 = n14002 & ~n14653;
  assign n15689 = ~n15687 & ~n15688;
  assign n15690 = n15686 & n15689;
  assign n15691 = n15683 & n15690;
  assign n15692 = n15676 & n15691;
  assign n15693 = n15671 & n15692;
  assign n15694 = ~n15657 & ~n15693;
  assign n15695 = n15618 & n15694;
  assign n15696 = ~n15546 & n15695;
  assign n15697 = pi021 & ~n11168;
  assign n15698 = n11073 & ~n11103;
  assign n15699 = n15697 & n15698;
  assign n15700 = ~n11188 & n15699;
  assign n15701 = ~n15620 & n15700;
  assign n15702 = ~n15619 & n15701;
  assign n15703 = ~n12380 & n15702;
  assign n15704 = ~n14467 & n15703;
  assign n15705 = ~n14466 & n15704;
  assign n15706 = n14574 & n15705;
  assign n15707 = n15629 & n15706;
  assign n15708 = n15633 & n15707;
  assign n15709 = n15595 & n15708;
  assign n15710 = n15656 & n15709;
  assign n15711 = pi023 & ~n12841;
  assign n15712 = n12775 & n15711;
  assign n15713 = ~n12902 & n15712;
  assign n15714 = ~n15659 & n15713;
  assign n15715 = ~n15658 & n15714;
  assign n15716 = ~n14467 & n15715;
  assign n15717 = ~n14466 & n15716;
  assign n15718 = n14574 & n15717;
  assign n15719 = n15666 & n15718;
  assign n15720 = n15669 & n15719;
  assign n15721 = n15595 & n15720;
  assign n15722 = n15692 & n15721;
  assign n15723 = ~n11551 & n14084;
  assign n15724 = ~n14467 & n15723;
  assign n15725 = ~n13906 & n15724;
  assign n15726 = ~n14452 & n15725;
  assign n15727 = n14456 & n15726;
  assign n15728 = n15571 & n15727;
  assign n15729 = n15585 & n15728;
  assign n15730 = ~n12471 & n12487;
  assign n15731 = ~n14467 & n15730;
  assign n15732 = ~n14466 & n15731;
  assign n15733 = n14574 & n15732;
  assign n15734 = n15599 & n15733;
  assign n15735 = n15595 & n15734;
  assign n15736 = n15593 & n15735;
  assign n15737 = n15615 & n15736;
  assign n15738 = ~n15729 & ~n15737;
  assign n15739 = ~n15722 & n15738;
  assign n15740 = ~n15710 & n15739;
  assign n15741 = ~n15696 & n15740;
  assign n15742 = n14382 & ~n14568;
  assign n15743 = ~n14320 & ~n14416;
  assign n15744 = ~n14350 & ~n14381;
  assign n15745 = n15743 & n15744;
  assign n15746 = ~n14519 & n15745;
  assign n15747 = ~n15742 & n15746;
  assign n15748 = ~n14467 & n15747;
  assign n15749 = ~n14466 & n15748;
  assign n15750 = n14574 & n15749;
  assign n15751 = ~n14577 & n15750;
  assign n15752 = ~n9717 & ~n9929;
  assign n15753 = ~n11266 & n15752;
  assign n15754 = ~n11588 & n15753;
  assign n15755 = ~n13859 & n15754;
  assign n15756 = ~n14676 & ~n15755;
  assign n15757 = n15751 & n15756;
  assign n15758 = n14457 & n15757;
  assign n15759 = ~n718 & ~n1372;
  assign n15760 = ~n2243 & n15759;
  assign n15761 = ~n3104 & n15760;
  assign n15762 = ~n3971 & n15761;
  assign n15763 = ~n4872 & n15762;
  assign n15764 = ~n5801 & n15763;
  assign n15765 = ~n6739 & n15764;
  assign n15766 = ~n7807 & n15765;
  assign n15767 = ~n8989 & n15766;
  assign n15768 = ~n10273 & n15767;
  assign n15769 = ~n11499 & n15768;
  assign n15770 = ~n13076 & n15769;
  assign n15771 = ~n14698 & n15770;
  assign n15772 = ~n6613 & ~n6784;
  assign n15773 = ~n7158 & n15772;
  assign n15774 = ~n8250 & n15773;
  assign n15775 = ~n9414 & n15774;
  assign n15776 = ~n10667 & n15775;
  assign n15777 = ~n12083 & n15776;
  assign n15778 = ~n13644 & n15777;
  assign n15779 = ~n10909 & ~n11188;
  assign n15780 = ~n12380 & n15779;
  assign n15781 = ~n14045 & n15780;
  assign n15782 = ~n15778 & ~n15781;
  assign n15783 = ~n15771 & n15782;
  assign n15784 = ~n5408 & ~n5808;
  assign n15785 = ~n6056 & n15784;
  assign n15786 = ~n7073 & n15785;
  assign n15787 = ~n8179 & n15786;
  assign n15788 = ~n9344 & n15787;
  assign n15789 = ~n10594 & n15788;
  assign n15790 = ~n12005 & n15789;
  assign n15791 = ~n13558 & n15790;
  assign n15792 = ~n4736 & ~n4817;
  assign n15793 = ~n4902 & n15792;
  assign n15794 = ~n6001 & n15793;
  assign n15795 = ~n7014 & n15794;
  assign n15796 = ~n8114 & n15795;
  assign n15797 = ~n9276 & n15796;
  assign n15798 = ~n10523 & n15797;
  assign n15799 = ~n11928 & n15798;
  assign n15800 = ~n13479 & n15799;
  assign n15801 = ~n15791 & ~n15800;
  assign n15802 = ~n3769 & ~n3940;
  assign n15803 = ~n4001 & n15802;
  assign n15804 = ~n5043 & n15803;
  assign n15805 = ~n5943 & n15804;
  assign n15806 = ~n6951 & n15805;
  assign n15807 = ~n8037 & n15806;
  assign n15808 = ~n9200 & n15807;
  assign n15809 = ~n10445 & n15808;
  assign n15810 = ~n11846 & n15809;
  assign n15811 = ~n13393 & n15810;
  assign n15812 = ~n1710 & ~n2242;
  assign n15813 = ~n3095 & n15812;
  assign n15814 = ~n3997 & n15813;
  assign n15815 = ~n4837 & n15814;
  assign n15816 = ~n5822 & n15815;
  assign n15817 = ~n6820 & n15816;
  assign n15818 = ~n7785 & n15817;
  assign n15819 = ~n9027 & n15818;
  assign n15820 = ~n10245 & n15819;
  assign n15821 = ~n11536 & n15820;
  assign n15822 = ~n13036 & n15821;
  assign n15823 = ~n14653 & n15822;
  assign n15824 = ~n15811 & ~n15823;
  assign n15825 = n15801 & n15824;
  assign n15826 = ~n12671 & ~n12902;
  assign n15827 = ~n14009 & n15826;
  assign n15828 = ~n7722 & ~n7869;
  assign n15829 = ~n8346 & n15828;
  assign n15830 = ~n9485 & n15829;
  assign n15831 = ~n10741 & n15830;
  assign n15832 = ~n12158 & n15831;
  assign n15833 = ~n13693 & n15832;
  assign n15834 = ~n15827 & ~n15833;
  assign n15835 = ~n2631 & ~n3066;
  assign n15836 = ~n3983 & n15835;
  assign n15837 = ~n4024 & n15836;
  assign n15838 = ~n4999 & n15837;
  assign n15839 = ~n5827 & n15838;
  assign n15840 = ~n6893 & n15839;
  assign n15841 = ~n7890 & n15840;
  assign n15842 = ~n9131 & n15841;
  assign n15843 = ~n10278 & n15842;
  assign n15844 = ~n11662 & n15843;
  assign n15845 = ~n13191 & n15844;
  assign n15846 = ~n8514 & ~n8834;
  assign n15847 = ~n10002 & n15846;
  assign n15848 = ~n11297 & n15847;
  assign n15849 = ~n12240 & n15848;
  assign n15850 = ~n13135 & n15849;
  assign n15851 = ~n15845 & ~n15850;
  assign n15852 = n15834 & n15851;
  assign n15853 = n15825 & n15852;
  assign n15854 = n15783 & n15853;
  assign n15855 = n15758 & n15854;
  assign n15856 = ~n12946 & ~n14467;
  assign n15857 = ~n14466 & n15856;
  assign n15858 = n14574 & n15857;
  assign n15859 = ~n13093 & ~n14451;
  assign n15860 = n15858 & n15859;
  assign n15861 = n12903 & ~n14009;
  assign n15862 = ~n14577 & ~n15861;
  assign n15863 = n15860 & n15862;
  assign n15864 = n15595 & n15863;
  assign n15865 = n12962 & ~n13393;
  assign n15866 = n13014 & ~n13644;
  assign n15867 = n13049 & ~n14045;
  assign n15868 = ~n15866 & ~n15867;
  assign n15869 = ~n15865 & n15868;
  assign n15870 = n13047 & ~n14653;
  assign n15871 = n12994 & ~n13135;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = n12986 & ~n13191;
  assign n15874 = n13088 & ~n14698;
  assign n15875 = ~n15873 & ~n15874;
  assign n15876 = n15872 & n15875;
  assign n15877 = n12970 & ~n13479;
  assign n15878 = n13008 & ~n13558;
  assign n15879 = ~n15877 & ~n15878;
  assign n15880 = n12989 & ~n13859;
  assign n15881 = n12999 & ~n13693;
  assign n15882 = ~n15880 & ~n15881;
  assign n15883 = n15879 & n15882;
  assign n15884 = n15876 & n15883;
  assign n15885 = n15869 & n15884;
  assign n15886 = n15864 & n15885;
  assign n15887 = ~n15855 & ~n15886;
  assign n15888 = ~n15741 & n15887;
  assign n15889 = pi025 & ~n14416;
  assign n15890 = n14351 & ~n14381;
  assign n15891 = n15889 & n15890;
  assign n15892 = ~n14519 & n15891;
  assign n15893 = ~n15742 & n15892;
  assign n15894 = ~n14467 & n15893;
  assign n15895 = ~n14466 & n15894;
  assign n15896 = n14574 & n15895;
  assign n15897 = ~n14577 & n15896;
  assign n15898 = n15756 & n15897;
  assign n15899 = n14457 & n15898;
  assign n15900 = n15854 & n15899;
  assign n15901 = n14118 & ~n14467;
  assign n15902 = ~n14466 & n15901;
  assign n15903 = n14574 & n15902;
  assign n15904 = n15859 & n15903;
  assign n15905 = n15862 & n15904;
  assign n15906 = n15595 & n15905;
  assign n15907 = n15885 & n15906;
  assign n15908 = ~n15900 & ~n15907;
  assign n15909 = ~n15888 & n15908;
  assign n15910 = ~n14716 & ~n15909;
  assign n15911 = pi026 & ~n14568;
  assign n15912 = ~n14520 & n15911;
  assign n15913 = ~n14467 & n15912;
  assign n15914 = ~n14466 & n15913;
  assign n15915 = n14574 & n15914;
  assign n15916 = ~n14465 & n15915;
  assign n15917 = n14581 & n15916;
  assign n15918 = n14457 & n15917;
  assign n15919 = n14715 & n15918;
  assign n15920 = n9854 & n11072;
  assign n15921 = n14178 & n15920;
  assign n15922 = ~pi249 & pi257;
  assign n15923 = pi249 & ~pi257;
  assign n15924 = ~pi250 & pi258;
  assign n15925 = pi250 & ~pi258;
  assign n15926 = ~pi251 & pi259;
  assign n15927 = pi251 & ~pi259;
  assign n15928 = ~pi252 & pi260;
  assign n15929 = pi252 & ~pi260;
  assign n15930 = pi254 & ~pi262;
  assign n15931 = pi253 & ~pi261;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = ~pi253 & pi261;
  assign n15934 = ~n15932 & ~n15933;
  assign n15935 = ~n15929 & ~n15934;
  assign n15936 = ~n15928 & ~n15935;
  assign n15937 = ~n15927 & ~n15936;
  assign n15938 = ~n15926 & ~n15937;
  assign n15939 = ~n15925 & ~n15938;
  assign n15940 = ~n15924 & ~n15939;
  assign n15941 = ~n15923 & ~n15940;
  assign n15942 = ~n15922 & ~n15941;
  assign n15943 = ~pi248 & ~n15942;
  assign n15944 = ~pi256 & ~n15943;
  assign n15945 = pi247 & ~pi255;
  assign n15946 = pi248 & ~n15922;
  assign n15947 = ~n15941 & n15946;
  assign n15948 = ~n15945 & ~n15947;
  assign n15949 = ~n15944 & n15948;
  assign n15950 = ~n14176 & ~n14415;
  assign n15951 = ~n15949 & n15950;
  assign n15952 = n12713 & n12811;
  assign n15953 = n15951 & n15952;
  assign n15954 = n15921 & n15953;
  assign n15955 = ~n1678 & ~n9653;
  assign n15956 = n12495 & n15955;
  assign n15957 = ~n1432 & ~n1739;
  assign n15958 = n10820 & n15957;
  assign n15959 = n15956 & n15958;
  assign n15960 = n10969 & n12641;
  assign n15961 = n9622 & n10818;
  assign n15962 = n15960 & n15961;
  assign n15963 = n15959 & n15962;
  assign n15964 = ~n2396 & ~n2515;
  assign n15965 = n3810 & n15964;
  assign n15966 = ~n1650 & ~n1711;
  assign n15967 = n2308 & n15966;
  assign n15968 = n15965 & n15967;
  assign n15969 = ~n3375 & ~n3563;
  assign n15970 = n14536 & n15969;
  assign n15971 = n14475 & n15970;
  assign n15972 = n15968 & n15971;
  assign n15973 = n12554 & n14521;
  assign n15974 = pi028 & ~n501;
  assign n15975 = n12872 & n15974;
  assign n15976 = n15973 & n15975;
  assign n15977 = n12559 & n12562;
  assign n15978 = ~n1209 & ~n2114;
  assign n15979 = n2311 & n15978;
  assign n15980 = n15977 & n15979;
  assign n15981 = n15976 & n15980;
  assign n15982 = n15972 & n15981;
  assign n15983 = ~n6314 & ~n7664;
  assign n15984 = n12545 & n15983;
  assign n15985 = ~n6465 & ~n6615;
  assign n15986 = n14201 & n15985;
  assign n15987 = n15984 & n15986;
  assign n15988 = ~n8456 & ~n14204;
  assign n15989 = ~pi247 & pi255;
  assign n15990 = ~n14387 & ~n15989;
  assign n15991 = n15988 & n15990;
  assign n15992 = n11400 & n14205;
  assign n15993 = n15991 & n15992;
  assign n15994 = n15987 & n15993;
  assign n15995 = ~n4283 & ~n4402;
  assign n15996 = ~n4679 & ~n5570;
  assign n15997 = n15995 & n15996;
  assign n15998 = ~n3256 & ~n3285;
  assign n15999 = n4796 & n15998;
  assign n16000 = n15997 & n15999;
  assign n16001 = ~n5350 & ~n5599;
  assign n16002 = n10836 & n16001;
  assign n16003 = n7242 & n16002;
  assign n16004 = n16000 & n16003;
  assign n16005 = n15994 & n16004;
  assign n16006 = n15982 & n16005;
  assign n16007 = ~n1172 & n16006;
  assign n16008 = ~n996 & n16007;
  assign n16009 = ~n2306 & n16008;
  assign n16010 = ~n500 & n16009;
  assign n16011 = ~n810 & ~n1237;
  assign n16012 = n16010 & n16011;
  assign n16013 = n12571 & n14143;
  assign n16014 = n6677 & n16013;
  assign n16015 = n16012 & n16014;
  assign n16016 = n10855 & n14185;
  assign n16017 = n14228 & n16016;
  assign n16018 = n16015 & n16017;
  assign n16019 = ~n6642 & ~n7691;
  assign n16020 = n14128 & n16019;
  assign n16021 = n10827 & n16020;
  assign n16022 = ~n8483 & ~n8542;
  assign n16023 = n12537 & n16022;
  assign n16024 = n14133 & n16023;
  assign n16025 = n16021 & n16024;
  assign n16026 = ~n2511 & ~n2542;
  assign n16027 = n5732 & n16026;
  assign n16028 = ~n3372 & ~n3590;
  assign n16029 = ~n3402 & ~n3738;
  assign n16030 = n16028 & n16029;
  assign n16031 = n16027 & n16030;
  assign n16032 = ~n5288 & ~n5626;
  assign n16033 = n14144 & n16032;
  assign n16034 = ~n4429 & ~n4607;
  assign n16035 = n14141 & n16034;
  assign n16036 = n16033 & n16035;
  assign n16037 = n16031 & n16036;
  assign n16038 = n16025 & n16037;
  assign n16039 = n16018 & n16038;
  assign n16040 = n15963 & n16039;
  assign n16041 = n15954 & n16040;
  assign n16042 = ~n6131 & n16041;
  assign n16043 = ~n14176 & ~n14319;
  assign n16044 = n12841 & n16043;
  assign n16045 = n11133 & n12811;
  assign n16046 = n9824 & n11103;
  assign n16047 = n16045 & n16046;
  assign n16048 = n16044 & n16047;
  assign n16049 = ~n2511 & ~n2571;
  assign n16050 = n5732 & n16049;
  assign n16051 = ~n3372 & ~n3619;
  assign n16052 = n16029 & n16051;
  assign n16053 = n16050 & n16052;
  assign n16054 = n16014 & n16053;
  assign n16055 = ~n2396 & ~n2544;
  assign n16056 = n3810 & n16055;
  assign n16057 = ~n1558 & ~n1650;
  assign n16058 = n2308 & n16057;
  assign n16059 = n16056 & n16058;
  assign n16060 = ~n3375 & ~n3592;
  assign n16061 = n14536 & n16060;
  assign n16062 = n14475 & n16061;
  assign n16063 = n16059 & n16062;
  assign n16064 = pi027 & ~n501;
  assign n16065 = n12872 & n16064;
  assign n16066 = n15973 & n16065;
  assign n16067 = ~n721 & ~n2114;
  assign n16068 = n2311 & n16067;
  assign n16069 = n15977 & n16068;
  assign n16070 = n16066 & n16069;
  assign n16071 = n16063 & n16070;
  assign n16072 = ~n7328 & ~n7447;
  assign n16073 = n11399 & n16072;
  assign n16074 = ~n6465 & ~n6556;
  assign n16075 = n14201 & n16074;
  assign n16076 = n16073 & n16075;
  assign n16077 = ~n8546 & ~n14204;
  assign n16078 = ~n14291 & n16077;
  assign n16079 = n15992 & n16078;
  assign n16080 = n16076 & n16079;
  assign n16081 = ~n4283 & ~n4461;
  assign n16082 = n15996 & n16081;
  assign n16083 = n15999 & n16082;
  assign n16084 = ~n5350 & ~n5629;
  assign n16085 = n10836 & n16084;
  assign n16086 = n7242 & n16085;
  assign n16087 = n16083 & n16086;
  assign n16088 = n16080 & n16087;
  assign n16089 = n16071 & n16088;
  assign n16090 = ~n1172 & n16089;
  assign n16091 = ~n996 & n16090;
  assign n16092 = ~n2306 & n16091;
  assign n16093 = ~n500 & n16092;
  assign n16094 = ~n749 & ~n810;
  assign n16095 = n16093 & n16094;
  assign n16096 = n16016 & n16095;
  assign n16097 = n16054 & n16096;
  assign n16098 = ~n8542 & ~n8573;
  assign n16099 = n12537 & n16098;
  assign n16100 = ~n7355 & ~n7474;
  assign n16101 = n10824 & n16100;
  assign n16102 = n16099 & n16101;
  assign n16103 = n9793 & n16102;
  assign n16104 = ~n5288 & ~n5656;
  assign n16105 = n14144 & n16104;
  assign n16106 = ~n4488 & ~n4607;
  assign n16107 = n14141 & n16106;
  assign n16108 = n16105 & n16107;
  assign n16109 = ~n6583 & ~n7750;
  assign n16110 = n14128 & n16109;
  assign n16111 = n10827 & n16110;
  assign n16112 = n16108 & n16111;
  assign n16113 = n16103 & n16112;
  assign n16114 = n16097 & n16113;
  assign n16115 = ~pi247 & pi271;
  assign n16116 = ~pi249 & pi273;
  assign n16117 = pi249 & ~pi273;
  assign n16118 = ~pi250 & pi274;
  assign n16119 = pi250 & ~pi274;
  assign n16120 = ~pi251 & pi275;
  assign n16121 = pi251 & ~pi275;
  assign n16122 = ~pi252 & pi276;
  assign n16123 = pi252 & ~pi276;
  assign n16124 = pi254 & ~pi278;
  assign n16125 = pi253 & ~pi277;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~pi253 & pi277;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = ~n16123 & ~n16128;
  assign n16130 = ~n16122 & ~n16129;
  assign n16131 = ~n16121 & ~n16130;
  assign n16132 = ~n16120 & ~n16131;
  assign n16133 = ~n16119 & ~n16132;
  assign n16134 = ~n16118 & ~n16133;
  assign n16135 = ~n16117 & ~n16134;
  assign n16136 = ~n16116 & ~n16135;
  assign n16137 = ~pi248 & ~n16136;
  assign n16138 = ~pi272 & ~n16137;
  assign n16139 = pi247 & ~pi271;
  assign n16140 = pi248 & ~n16116;
  assign n16141 = ~n16135 & n16140;
  assign n16142 = ~n16139 & ~n16141;
  assign n16143 = ~n16138 & n16142;
  assign n16144 = ~n16115 & ~n16143;
  assign n16145 = n15960 & ~n16144;
  assign n16146 = ~pi247 & pi263;
  assign n16147 = ~pi249 & pi265;
  assign n16148 = pi249 & ~pi265;
  assign n16149 = ~pi250 & pi266;
  assign n16150 = pi250 & ~pi266;
  assign n16151 = ~pi251 & pi267;
  assign n16152 = pi251 & ~pi267;
  assign n16153 = ~pi252 & pi268;
  assign n16154 = pi252 & ~pi268;
  assign n16155 = pi254 & ~pi270;
  assign n16156 = pi253 & ~pi269;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = ~pi253 & pi269;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = ~n16154 & ~n16159;
  assign n16161 = ~n16153 & ~n16160;
  assign n16162 = ~n16152 & ~n16161;
  assign n16163 = ~n16151 & ~n16162;
  assign n16164 = ~n16150 & ~n16163;
  assign n16165 = ~n16149 & ~n16164;
  assign n16166 = ~n16148 & ~n16165;
  assign n16167 = ~n16147 & ~n16166;
  assign n16168 = ~pi248 & ~n16167;
  assign n16169 = ~pi264 & ~n16168;
  assign n16170 = pi247 & ~pi263;
  assign n16171 = pi248 & ~n16147;
  assign n16172 = ~n16166 & n16171;
  assign n16173 = ~n16170 & ~n16172;
  assign n16174 = ~n16169 & n16173;
  assign n16175 = ~n16146 & ~n16174;
  assign n16176 = ~n15949 & ~n15989;
  assign n16177 = ~n16175 & ~n16176;
  assign n16178 = n16145 & n16177;
  assign n16179 = ~n1432 & ~n1586;
  assign n16180 = n10820 & n16179;
  assign n16181 = n14228 & n16180;
  assign n16182 = n15956 & n15961;
  assign n16183 = n16181 & n16182;
  assign n16184 = n16178 & n16183;
  assign n16185 = n16114 & n16184;
  assign n16186 = n16048 & n16185;
  assign n16187 = ~n6131 & n16186;
  assign n16188 = ~n16042 & ~n16187;
  assign n16189 = ~n6137 & ~n7236;
  assign n16190 = ~n6125 & ~n6132;
  assign n16191 = n6193 & n16190;
  assign n16192 = n16189 & n16191;
  assign n16193 = ~n16188 & n16192;
  assign n16194 = ~n8867 & n16193;
  assign n16195 = ~n7235 & n16194;
  assign n16196 = n7296 & n16195;
  assign n16197 = n7231 & n16196;
  assign n16198 = ~n10027 & n16197;
  assign n16199 = ~n8866 & n16198;
  assign n16200 = n8898 & n16199;
  assign n16201 = n8863 & n16200;
  assign n16202 = ~n10788 & n16201;
  assign n16203 = ~n10026 & n16202;
  assign n16204 = n10072 & n16203;
  assign n16205 = n10021 & n16204;
  assign n16206 = ~n15919 & ~n16205;
  assign po014 = n15910 | ~n16206;
  assign n16208 = n14452 & ~n14741;
  assign n16209 = n14455 & ~n15419;
  assign n16210 = ~n16208 & ~n16209;
  assign n16211 = n14454 & ~n15465;
  assign n16212 = n14577 & ~n15616;
  assign n16213 = ~n16211 & ~n16212;
  assign n16214 = n16210 & n16213;
  assign n16215 = n14572 & ~n15167;
  assign n16216 = n14467 & ~n14980;
  assign n16217 = ~pi026 & ~n14568;
  assign n16218 = ~n16216 & n16217;
  assign n16219 = ~n16215 & n16218;
  assign n16220 = n14573 & ~n15075;
  assign n16221 = n14466 & ~n15278;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = n16219 & n16222;
  assign n16224 = n14451 & ~n15586;
  assign n16225 = ~n14716 & ~n16224;
  assign n16226 = n16223 & n16225;
  assign n16227 = n14625 & ~n14848;
  assign n16228 = n14580 & ~n15657;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = n16226 & n16229;
  assign n16231 = n16214 & n16230;
  assign n16232 = n14676 & ~n15886;
  assign n16233 = n14520 & ~n15855;
  assign n16234 = ~n16232 & ~n16233;
  assign n16235 = ~n2242 & n3070;
  assign n16236 = ~n3095 & n16235;
  assign n16237 = ~n3997 & n16236;
  assign n16238 = ~n4003 & n16237;
  assign n16239 = ~n4837 & n16238;
  assign n16240 = ~n5822 & n16239;
  assign n16241 = ~n6820 & n16240;
  assign n16242 = ~n7785 & n16241;
  assign n16243 = ~n9027 & n16242;
  assign n16244 = ~n10245 & n16243;
  assign n16245 = ~n14919 & n16244;
  assign n16246 = ~n14918 & n16245;
  assign n16247 = ~n11536 & n16246;
  assign n16248 = ~n13036 & n16247;
  assign n16249 = ~n14917 & n16248;
  assign n16250 = ~n14916 & n16249;
  assign n16251 = n14940 & n16250;
  assign n16252 = n14943 & n16251;
  assign n16253 = n14947 & n16252;
  assign n16254 = n14915 & n16253;
  assign n16255 = n14970 & n16254;
  assign n16256 = n14665 & ~n16255;
  assign n16257 = n14592 & ~n15153;
  assign n16258 = ~n16256 & ~n16257;
  assign n16259 = n16234 & n16258;
  assign n16260 = n14465 & ~n15239;
  assign n16261 = n14598 & ~n15385;
  assign n16262 = ~n16260 & ~n16261;
  assign n16263 = n14614 & ~n15061;
  assign n16264 = ~n1372 & n2272;
  assign n16265 = ~n2243 & n16264;
  assign n16266 = ~n3104 & n16265;
  assign n16267 = ~n3837 & n16266;
  assign n16268 = ~n3971 & n16267;
  assign n16269 = ~n4872 & n16268;
  assign n16270 = ~n5801 & n16269;
  assign n16271 = ~n6739 & n16270;
  assign n16272 = ~n7807 & n16271;
  assign n16273 = ~n8989 & n16272;
  assign n16274 = ~n10273 & n16273;
  assign n16275 = ~n14857 & n16274;
  assign n16276 = ~n14856 & n16275;
  assign n16277 = ~n11499 & n16276;
  assign n16278 = ~n13076 & n16277;
  assign n16279 = ~n14855 & n16278;
  assign n16280 = ~n14854 & n16279;
  assign n16281 = n14879 & n16280;
  assign n16282 = n14882 & n16281;
  assign n16283 = n14886 & n16282;
  assign n16284 = n14853 & n16283;
  assign n16285 = n14909 & n16284;
  assign n16286 = n14711 & ~n16285;
  assign n16287 = ~n16263 & ~n16286;
  assign n16288 = n16262 & n16287;
  assign n16289 = n14602 & ~n15536;
  assign n16290 = n14674 & ~n15693;
  assign n16291 = ~n16289 & ~n16290;
  assign n16292 = n14633 & ~n15330;
  assign n16293 = n14672 & ~n15482;
  assign n16294 = ~n16292 & ~n16293;
  assign n16295 = n16291 & n16294;
  assign n16296 = n16288 & n16295;
  assign n16297 = n16259 & n16296;
  assign n16298 = n16231 & n16297;
  assign n16299 = ~n14741 & n15189;
  assign n16300 = n15191 & ~n15419;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = n15210 & ~n15586;
  assign n16303 = n15223 & ~n15616;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = n16301 & n16304;
  assign n16306 = n3859 & n14194;
  assign n16307 = n12916 & n16057;
  assign n16308 = n16306 & n16307;
  assign n16309 = n7812 & n16061;
  assign n16310 = n16308 & n16309;
  assign n16311 = n10840 & n16067;
  assign n16312 = n2246 & n16311;
  assign n16313 = ~n504 & ~n659;
  assign n16314 = n12554 & n16313;
  assign n16315 = n5755 & n16314;
  assign n16316 = n16312 & n16315;
  assign n16317 = n16310 & n16316;
  assign n16318 = n8868 & n16072;
  assign n16319 = ~n6494 & ~n6556;
  assign n16320 = n12544 & n16319;
  assign n16321 = n16318 & n16320;
  assign n16322 = ~n8515 & ~n14291;
  assign n16323 = n16077 & n16322;
  assign n16324 = ~n7387 & ~n7723;
  assign n16325 = n12904 & n16324;
  assign n16326 = n16323 & n16325;
  assign n16327 = n16321 & n16326;
  assign n16328 = ~n2544 & ~n3227;
  assign n16329 = n14210 & n16328;
  assign n16330 = n16082 & n16329;
  assign n16331 = n6741 & n16085;
  assign n16332 = n16330 & n16331;
  assign n16333 = n16327 & n16332;
  assign n16334 = n16317 & n16333;
  assign n16335 = ~n1172 & n16334;
  assign n16336 = ~n996 & n16335;
  assign n16337 = ~n2306 & n16336;
  assign n16338 = ~n500 & n16337;
  assign n16339 = n16094 & n16338;
  assign n16340 = n16016 & n16339;
  assign n16341 = n16054 & n16340;
  assign n16342 = n16113 & n16341;
  assign n16343 = n16184 & n16342;
  assign n16344 = n16048 & n16343;
  assign n16345 = ~n7236 & n16344;
  assign n16346 = ~n6137 & n16345;
  assign n16347 = n6193 & n16346;
  assign n16348 = n6134 & n16347;
  assign n16349 = ~n8867 & n16348;
  assign n16350 = ~n7235 & n16349;
  assign n16351 = n7296 & n16350;
  assign n16352 = n7231 & n16351;
  assign n16353 = ~n10027 & n16352;
  assign n16354 = ~n8866 & n16353;
  assign n16355 = n8898 & n16354;
  assign n16356 = n8863 & n16355;
  assign n16357 = ~n10788 & n16356;
  assign n16358 = ~n10026 & n16357;
  assign n16359 = n10072 & n16358;
  assign n16360 = n10021 & n16359;
  assign n16361 = n5657 & ~n16360;
  assign n16362 = n3941 & n14194;
  assign n16363 = ~n2515 & ~n3227;
  assign n16364 = n12916 & n16363;
  assign n16365 = n16362 & n16364;
  assign n16366 = n14275 & n15970;
  assign n16367 = n16365 & n16366;
  assign n16368 = n10840 & n16313;
  assign n16369 = n2246 & n15978;
  assign n16370 = n16368 & n16369;
  assign n16371 = n5717 & n15966;
  assign n16372 = n5754 & n12554;
  assign n16373 = n16371 & n16372;
  assign n16374 = n16370 & n16373;
  assign n16375 = n16367 & n16374;
  assign n16376 = ~n7328 & ~n7723;
  assign n16377 = ~n7387 & ~n7664;
  assign n16378 = n16376 & n16377;
  assign n16379 = n8869 & n16378;
  assign n16380 = ~n8515 & ~n14387;
  assign n16381 = ~n15989 & n16380;
  assign n16382 = n12904 & n15988;
  assign n16383 = n16381 & n16382;
  assign n16384 = n16379 & n16383;
  assign n16385 = n12909 & n15997;
  assign n16386 = ~n6494 & ~n6615;
  assign n16387 = n16001 & n16386;
  assign n16388 = n12906 & n16387;
  assign n16389 = n16385 & n16388;
  assign n16390 = n16384 & n16389;
  assign n16391 = n16375 & n16390;
  assign n16392 = ~n1172 & n16391;
  assign n16393 = ~n996 & n16392;
  assign n16394 = ~n2306 & n16393;
  assign n16395 = ~n500 & n16394;
  assign n16396 = n16011 & n16395;
  assign n16397 = n16014 & n16396;
  assign n16398 = n16017 & n16397;
  assign n16399 = n16038 & n16398;
  assign n16400 = n15963 & n16399;
  assign n16401 = n15954 & n16400;
  assign n16402 = ~n7236 & n16401;
  assign n16403 = ~n6137 & n16402;
  assign n16404 = n6193 & n16403;
  assign n16405 = n6134 & n16404;
  assign n16406 = ~n8867 & n16405;
  assign n16407 = ~n7235 & n16406;
  assign n16408 = n7296 & n16407;
  assign n16409 = n7231 & n16408;
  assign n16410 = ~n10027 & n16409;
  assign n16411 = ~n8866 & n16410;
  assign n16412 = n8898 & n16411;
  assign n16413 = n8863 & n16412;
  assign n16414 = ~n10788 & n16413;
  assign n16415 = ~n10026 & n16414;
  assign n16416 = n10072 & n16415;
  assign n16417 = n10021 & n16416;
  assign n16418 = n5627 & ~n16417;
  assign n16419 = ~n5808 & n6064;
  assign n16420 = ~n6056 & n16419;
  assign n16421 = ~n7073 & n16420;
  assign n16422 = ~n8179 & n16421;
  assign n16423 = ~n9344 & n16422;
  assign n16424 = ~n16418 & n16423;
  assign n16425 = ~n16361 & n16424;
  assign n16426 = ~n10594 & n16425;
  assign n16427 = ~n12005 & n16426;
  assign n16428 = ~n13558 & n16427;
  assign n16429 = ~n16216 & n16428;
  assign n16430 = ~n16215 & n16429;
  assign n16431 = n15207 & ~n15278;
  assign n16432 = ~n16220 & ~n16431;
  assign n16433 = n16430 & n16432;
  assign n16434 = n15190 & ~n15465;
  assign n16435 = ~n15239 & ~n16434;
  assign n16436 = n16433 & n16435;
  assign n16437 = n15218 & ~n15886;
  assign n16438 = n15194 & ~n15855;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = n16436 & n16439;
  assign n16441 = n16305 & n16440;
  assign n16442 = n15220 & ~n16285;
  assign n16443 = ~n14848 & n15233;
  assign n16444 = ~n16442 & ~n16443;
  assign n16445 = ~n15061 & n15219;
  assign n16446 = n15230 & ~n15482;
  assign n16447 = ~n16445 & ~n16446;
  assign n16448 = n16444 & n16447;
  assign n16449 = ~n14716 & n15195;
  assign n16450 = n15224 & ~n15385;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = n15226 & ~n15657;
  assign n16453 = n15213 & ~n15536;
  assign n16454 = ~n16452 & ~n16453;
  assign n16455 = n16451 & n16454;
  assign n16456 = ~n15153 & n15234;
  assign n16457 = n15231 & ~n15693;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = n15214 & ~n16255;
  assign n16460 = n15227 & ~n15330;
  assign n16461 = ~n16459 & ~n16460;
  assign n16462 = n16458 & n16461;
  assign n16463 = n16455 & n16462;
  assign n16464 = n16448 & n16463;
  assign n16465 = n16441 & n16464;
  assign n16466 = n15160 & ~n16285;
  assign n16467 = n16215 & ~n16216;
  assign n16468 = ~n16220 & n16467;
  assign n16469 = ~n16466 & n16468;
  assign n16470 = ~n14848 & n15164;
  assign n16471 = ~n15061 & n15163;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = n15156 & ~n16255;
  assign n16474 = ~n15153 & n15161;
  assign n16475 = ~n16473 & ~n16474;
  assign n16476 = n16472 & n16475;
  assign n16477 = n16469 & n16476;
  assign n16478 = ~n14741 & n15102;
  assign n16479 = n15101 & ~n15465;
  assign n16480 = ~n16478 & ~n16479;
  assign n16481 = n15124 & ~n15586;
  assign n16482 = n15127 & ~n15616;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = n16480 & n16483;
  assign n16485 = n4430 & ~n16417;
  assign n16486 = n4489 & ~n16360;
  assign n16487 = ~n4401 & ~n4460;
  assign n16488 = ~n4817 & n16487;
  assign n16489 = ~n4902 & n16488;
  assign n16490 = ~n6001 & n16489;
  assign n16491 = ~n7014 & n16490;
  assign n16492 = ~n8114 & n16491;
  assign n16493 = ~n9276 & n16492;
  assign n16494 = ~n16486 & n16493;
  assign n16495 = ~n16485 & n16494;
  assign n16496 = ~n10523 & n16495;
  assign n16497 = ~n11928 & n16496;
  assign n16498 = ~n13479 & n16497;
  assign n16499 = ~n16216 & n16498;
  assign n16500 = ~n16220 & n16499;
  assign n16501 = n15120 & ~n15167;
  assign n16502 = n15121 & ~n15278;
  assign n16503 = ~n16501 & ~n16502;
  assign n16504 = n16500 & n16503;
  assign n16505 = n15103 & ~n15419;
  assign n16506 = ~n15153 & ~n16505;
  assign n16507 = n16504 & n16506;
  assign n16508 = n15132 & ~n15886;
  assign n16509 = n15106 & ~n15855;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = n16507 & n16510;
  assign n16512 = n16484 & n16511;
  assign n16513 = n15134 & ~n16285;
  assign n16514 = ~n14848 & n15141;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = ~n15061 & n15138;
  assign n16517 = n15148 & ~n15482;
  assign n16518 = ~n16516 & ~n16517;
  assign n16519 = n16515 & n16518;
  assign n16520 = ~n14716 & n15107;
  assign n16521 = n15128 & ~n15385;
  assign n16522 = ~n16520 & ~n16521;
  assign n16523 = n15140 & ~n15657;
  assign n16524 = n15137 & ~n15536;
  assign n16525 = ~n16523 & ~n16524;
  assign n16526 = n16522 & n16525;
  assign n16527 = n15133 & ~n15239;
  assign n16528 = n15145 & ~n15693;
  assign n16529 = ~n16527 & ~n16528;
  assign n16530 = n15144 & ~n16255;
  assign n16531 = n15147 & ~n15330;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = n16529 & n16532;
  assign n16534 = n16526 & n16533;
  assign n16535 = n16519 & n16534;
  assign n16536 = n16512 & n16535;
  assign n16537 = ~n15061 & n15071;
  assign n16538 = ~n16216 & n16220;
  assign n16539 = ~n16537 & n16538;
  assign n16540 = n15070 & ~n16285;
  assign n16541 = ~n14848 & n15072;
  assign n16542 = n15067 & ~n16255;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = ~n16540 & n16543;
  assign n16545 = n16539 & n16544;
  assign n16546 = ~n14741 & n15007;
  assign n16547 = n15006 & ~n15465;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = n15005 & ~n15419;
  assign n16550 = n15032 & ~n15586;
  assign n16551 = ~n16549 & ~n16550;
  assign n16552 = n16548 & n16551;
  assign n16553 = n15028 & ~n15167;
  assign n16554 = n3620 & ~n16360;
  assign n16555 = n3591 & ~n16417;
  assign n16556 = ~n3650 & n10461;
  assign n16557 = ~n3940 & n16556;
  assign n16558 = ~n4001 & n16557;
  assign n16559 = ~n5043 & n16558;
  assign n16560 = ~n5943 & n16559;
  assign n16561 = ~n6951 & n16560;
  assign n16562 = ~n8037 & n16561;
  assign n16563 = ~n9200 & n16562;
  assign n16564 = ~n16555 & n16563;
  assign n16565 = ~n16554 & n16564;
  assign n16566 = ~n10445 & n16565;
  assign n16567 = ~n11846 & n16566;
  assign n16568 = ~n13393 & n16567;
  assign n16569 = ~n16216 & n16568;
  assign n16570 = ~n16553 & n16569;
  assign n16571 = n15010 & ~n15075;
  assign n16572 = n15029 & ~n15278;
  assign n16573 = ~n16571 & ~n16572;
  assign n16574 = n16570 & n16573;
  assign n16575 = n15053 & ~n15616;
  assign n16576 = ~n15061 & ~n16575;
  assign n16577 = n16574 & n16576;
  assign n16578 = ~n14716 & n15011;
  assign n16579 = n15012 & ~n15855;
  assign n16580 = ~n16578 & ~n16579;
  assign n16581 = n16577 & n16580;
  assign n16582 = n16552 & n16581;
  assign n16583 = n15045 & ~n16255;
  assign n16584 = ~n14848 & n15041;
  assign n16585 = ~n16583 & ~n16584;
  assign n16586 = n15046 & ~n15239;
  assign n16587 = n15035 & ~n15153;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = n16585 & n16588;
  assign n16590 = n15042 & ~n16285;
  assign n16591 = n15049 & ~n15330;
  assign n16592 = ~n16590 & ~n16591;
  assign n16593 = n15055 & ~n15536;
  assign n16594 = n15048 & ~n15657;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = n16592 & n16595;
  assign n16597 = n15040 & ~n15886;
  assign n16598 = n15052 & ~n15482;
  assign n16599 = ~n16597 & ~n16598;
  assign n16600 = n15036 & ~n15385;
  assign n16601 = n15056 & ~n15693;
  assign n16602 = ~n16600 & ~n16601;
  assign n16603 = n16599 & n16602;
  assign n16604 = n16596 & n16603;
  assign n16605 = n16589 & n16604;
  assign n16606 = n16582 & n16605;
  assign n16607 = n14791 & ~n15419;
  assign n16608 = n14790 & ~n15465;
  assign n16609 = ~n16607 & ~n16608;
  assign n16610 = ~n14741 & n14789;
  assign n16611 = n14832 & ~n15616;
  assign n16612 = ~n16610 & ~n16611;
  assign n16613 = n16609 & n16612;
  assign n16614 = n14794 & ~n15075;
  assign n16615 = n14795 & ~n14980;
  assign n16616 = n2543 & ~n16417;
  assign n16617 = n2572 & ~n16360;
  assign n16618 = ~n3066 & n14798;
  assign n16619 = ~n3983 & n16618;
  assign n16620 = ~n4003 & n16619;
  assign n16621 = ~n4024 & n16620;
  assign n16622 = ~n4999 & n16621;
  assign n16623 = ~n5827 & n16622;
  assign n16624 = ~n6893 & n16623;
  assign n16625 = ~n7890 & n16624;
  assign n16626 = ~n9131 & n16625;
  assign n16627 = ~n16617 & n16626;
  assign n16628 = ~n16616 & n16627;
  assign n16629 = ~n10278 & n16628;
  assign n16630 = ~n11662 & n16629;
  assign n16631 = ~n13191 & n16630;
  assign n16632 = ~n16615 & n16631;
  assign n16633 = ~n16614 & n16632;
  assign n16634 = n14816 & ~n15278;
  assign n16635 = n14815 & ~n15167;
  assign n16636 = ~n16634 & ~n16635;
  assign n16637 = n16633 & n16636;
  assign n16638 = n14819 & ~n15586;
  assign n16639 = ~n14848 & ~n16638;
  assign n16640 = n16637 & n16639;
  assign n16641 = n14796 & ~n15855;
  assign n16642 = ~n14716 & n14797;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = n16640 & n16643;
  assign n16645 = n16613 & n16644;
  assign n16646 = n14839 & ~n15482;
  assign n16647 = n14840 & ~n15153;
  assign n16648 = ~n16646 & ~n16647;
  assign n16649 = n14843 & ~n15061;
  assign n16650 = n14828 & ~n15536;
  assign n16651 = ~n16649 & ~n16650;
  assign n16652 = n16648 & n16651;
  assign n16653 = n14822 & ~n16255;
  assign n16654 = n14823 & ~n15693;
  assign n16655 = ~n16653 & ~n16654;
  assign n16656 = n14836 & ~n15239;
  assign n16657 = n14833 & ~n15385;
  assign n16658 = ~n16656 & ~n16657;
  assign n16659 = n16655 & n16658;
  assign n16660 = n14835 & ~n15657;
  assign n16661 = n14842 & ~n15330;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = n14829 & ~n16285;
  assign n16664 = n14827 & ~n15886;
  assign n16665 = ~n16663 & ~n16664;
  assign n16666 = n16662 & n16665;
  assign n16667 = n16659 & n16666;
  assign n16668 = n16652 & n16667;
  assign n16669 = n16645 & n16668;
  assign n16670 = n14881 & ~n15586;
  assign n16671 = n14851 & ~n15465;
  assign n16672 = ~n16670 & ~n16671;
  assign n16673 = ~n14741 & n14850;
  assign n16674 = n14849 & ~n15419;
  assign n16675 = ~n16673 & ~n16674;
  assign n16676 = n16672 & n16675;
  assign n16677 = n14877 & ~n15278;
  assign n16678 = n14855 & ~n14980;
  assign n16679 = n750 & ~n16360;
  assign n16680 = n1238 & ~n16417;
  assign n16681 = n2264 & ~n3828;
  assign n16682 = ~n4002 & n16681;
  assign n16683 = ~n780 & n10294;
  assign n16684 = ~n1372 & n16683;
  assign n16685 = ~n2243 & n16684;
  assign n16686 = ~n3104 & n16685;
  assign n16687 = ~n3971 & n16686;
  assign n16688 = ~n16682 & n16687;
  assign n16689 = ~n4872 & n16688;
  assign n16690 = ~n5801 & n16689;
  assign n16691 = ~n6739 & n16690;
  assign n16692 = ~n7807 & n16691;
  assign n16693 = ~n8989 & n16692;
  assign n16694 = ~n10273 & n16693;
  assign n16695 = ~n16680 & n16694;
  assign n16696 = ~n16679 & n16695;
  assign n16697 = ~n11499 & n16696;
  assign n16698 = ~n13076 & n16697;
  assign n16699 = ~n14698 & n16698;
  assign n16700 = ~n16678 & n16699;
  assign n16701 = ~n16677 & n16700;
  assign n16702 = n14854 & ~n15167;
  assign n16703 = n14878 & ~n15075;
  assign n16704 = ~n16702 & ~n16703;
  assign n16705 = n16701 & n16704;
  assign n16706 = n14884 & ~n15616;
  assign n16707 = ~n16285 & ~n16706;
  assign n16708 = n16705 & n16707;
  assign n16709 = n14889 & ~n15886;
  assign n16710 = n14894 & ~n15061;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = n16708 & n16711;
  assign n16713 = n16676 & n16712;
  assign n16714 = n14901 & ~n15330;
  assign n16715 = n14902 & ~n15536;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = n14857 & ~n15855;
  assign n16718 = ~n14716 & n14856;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = n16716 & n16719;
  assign n16721 = n14897 & ~n15657;
  assign n16722 = n14891 & ~n15693;
  assign n16723 = ~n16721 & ~n16722;
  assign n16724 = n14905 & ~n15239;
  assign n16725 = n14898 & ~n15385;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = n16723 & n16726;
  assign n16728 = n14885 & ~n15153;
  assign n16729 = ~n14848 & n14895;
  assign n16730 = ~n16728 & ~n16729;
  assign n16731 = n14904 & ~n15482;
  assign n16732 = n14890 & ~n16255;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = n16730 & n16733;
  assign n16735 = n16727 & n16734;
  assign n16736 = n16720 & n16735;
  assign n16737 = n16713 & n16736;
  assign n16738 = n14913 & ~n15465;
  assign n16739 = ~n14741 & n14942;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = n14912 & ~n15586;
  assign n16742 = n14963 & ~n15616;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 = n16740 & n16743;
  assign n16745 = n14938 & ~n15075;
  assign n16746 = n14917 & ~n14980;
  assign n16747 = n1587 & ~n16360;
  assign n16748 = n1740 & ~n16417;
  assign n16749 = pi003 & ~n1526;
  assign n16750 = ~n1556 & n16749;
  assign n16751 = ~n2242 & n16750;
  assign n16752 = ~n3095 & n16751;
  assign n16753 = ~n3997 & n16752;
  assign n16754 = ~n4003 & n16753;
  assign n16755 = ~n4837 & n16754;
  assign n16756 = ~n5822 & n16755;
  assign n16757 = ~n6820 & n16756;
  assign n16758 = ~n7785 & n16757;
  assign n16759 = ~n9027 & n16758;
  assign n16760 = ~n10245 & n16759;
  assign n16761 = ~n16748 & n16760;
  assign n16762 = ~n16747 & n16761;
  assign n16763 = ~n11536 & n16762;
  assign n16764 = ~n13036 & n16763;
  assign n16765 = ~n14653 & n16764;
  assign n16766 = ~n16746 & n16765;
  assign n16767 = ~n16745 & n16766;
  assign n16768 = n14916 & ~n15278;
  assign n16769 = n14939 & ~n15167;
  assign n16770 = ~n16768 & ~n16769;
  assign n16771 = n16767 & n16770;
  assign n16772 = n14911 & ~n15419;
  assign n16773 = ~n16255 & ~n16772;
  assign n16774 = n16771 & n16773;
  assign n16775 = ~n14848 & n14966;
  assign n16776 = n14956 & ~n15061;
  assign n16777 = ~n16775 & ~n16776;
  assign n16778 = n16774 & n16777;
  assign n16779 = n16744 & n16778;
  assign n16780 = n14951 & ~n15385;
  assign n16781 = n14946 & ~n15330;
  assign n16782 = ~n16780 & ~n16781;
  assign n16783 = n14919 & ~n15855;
  assign n16784 = ~n14716 & n14918;
  assign n16785 = ~n16783 & ~n16784;
  assign n16786 = n16782 & n16785;
  assign n16787 = n14962 & ~n15693;
  assign n16788 = n14958 & ~n15657;
  assign n16789 = ~n16787 & ~n16788;
  assign n16790 = n14945 & ~n15536;
  assign n16791 = n14955 & ~n15482;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = n16789 & n16792;
  assign n16794 = n14959 & ~n15239;
  assign n16795 = n14965 & ~n15153;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = n14952 & ~n16285;
  assign n16798 = n14950 & ~n15886;
  assign n16799 = ~n16797 & ~n16798;
  assign n16800 = n16796 & n16799;
  assign n16801 = n16793 & n16800;
  assign n16802 = n16786 & n16801;
  assign n16803 = n16779 & n16802;
  assign n16804 = ~n16737 & ~n16803;
  assign n16805 = ~n16669 & n16804;
  assign n16806 = ~pi005 & ~n2602;
  assign n16807 = ~n2783 & n16806;
  assign n16808 = ~n3066 & n16807;
  assign n16809 = ~n3983 & n16808;
  assign n16810 = ~n4003 & n16809;
  assign n16811 = ~n4024 & n16810;
  assign n16812 = ~n4999 & n16811;
  assign n16813 = ~n5827 & n16812;
  assign n16814 = ~n6893 & n16813;
  assign n16815 = ~n7890 & n16814;
  assign n16816 = ~n9131 & n16815;
  assign n16817 = ~n16617 & n16816;
  assign n16818 = ~n16616 & n16817;
  assign n16819 = ~n10278 & n16818;
  assign n16820 = ~n11662 & n16819;
  assign n16821 = ~n13191 & n16820;
  assign n16822 = ~n16615 & n16821;
  assign n16823 = ~n16614 & n16822;
  assign n16824 = n16636 & n16823;
  assign n16825 = n16639 & n16824;
  assign n16826 = n16643 & n16825;
  assign n16827 = n16613 & n16826;
  assign n16828 = n16668 & n16827;
  assign n16829 = n14978 & ~n16255;
  assign n16830 = ~n14974 & ~n14977;
  assign n16831 = ~n14978 & n16830;
  assign n16832 = n14975 & ~n16831;
  assign n16833 = ~n16829 & n16832;
  assign n16834 = ~n14848 & n14977;
  assign n16835 = n14974 & ~n16285;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = n16833 & n16836;
  assign n16838 = ~n16828 & ~n16837;
  assign n16839 = ~n16805 & n16838;
  assign n16840 = ~n3650 & ~n3710;
  assign n16841 = ~n3940 & n16840;
  assign n16842 = ~n4001 & n16841;
  assign n16843 = ~n5043 & n16842;
  assign n16844 = ~n5943 & n16843;
  assign n16845 = ~n6951 & n16844;
  assign n16846 = ~n8037 & n16845;
  assign n16847 = ~n9200 & n16846;
  assign n16848 = ~n16555 & n16847;
  assign n16849 = ~n16554 & n16848;
  assign n16850 = ~n10445 & n16849;
  assign n16851 = ~n11846 & n16850;
  assign n16852 = ~n13393 & n16851;
  assign n16853 = ~n16216 & n16852;
  assign n16854 = ~n16553 & n16853;
  assign n16855 = n16573 & n16854;
  assign n16856 = n16576 & n16855;
  assign n16857 = n16580 & n16856;
  assign n16858 = n16552 & n16857;
  assign n16859 = n16605 & n16858;
  assign n16860 = n15062 & ~n16831;
  assign n16861 = ~n16829 & n16860;
  assign n16862 = n16836 & n16861;
  assign n16863 = ~n16859 & ~n16862;
  assign n16864 = ~n16839 & n16863;
  assign n16865 = ~n16606 & ~n16864;
  assign n16866 = ~n16545 & ~n16865;
  assign n16867 = ~n6967 & n6983;
  assign n16868 = ~n8053 & n16867;
  assign n16869 = ~n9215 & n16868;
  assign n16870 = ~n10460 & n16869;
  assign n16871 = ~n11860 & n16870;
  assign n16872 = ~n13407 & n16871;
  assign n16873 = ~n15075 & n16872;
  assign n16874 = ~n16216 & n16873;
  assign n16875 = ~n16537 & n16874;
  assign n16876 = n16544 & n16875;
  assign n16877 = ~n16866 & ~n16876;
  assign n16878 = ~n16536 & ~n16877;
  assign n16879 = ~n4460 & n15168;
  assign n16880 = ~n4817 & n16879;
  assign n16881 = ~n4902 & n16880;
  assign n16882 = ~n6001 & n16881;
  assign n16883 = ~n7014 & n16882;
  assign n16884 = ~n8114 & n16883;
  assign n16885 = ~n9276 & n16884;
  assign n16886 = ~n16486 & n16885;
  assign n16887 = ~n16485 & n16886;
  assign n16888 = ~n10523 & n16887;
  assign n16889 = ~n11928 & n16888;
  assign n16890 = ~n13479 & n16889;
  assign n16891 = ~n16216 & n16890;
  assign n16892 = ~n16220 & n16891;
  assign n16893 = n16503 & n16892;
  assign n16894 = n16506 & n16893;
  assign n16895 = n16510 & n16894;
  assign n16896 = n16484 & n16895;
  assign n16897 = n16535 & n16896;
  assign n16898 = ~n16878 & ~n16897;
  assign n16899 = ~n16477 & ~n16898;
  assign n16900 = ~n7029 & n7074;
  assign n16901 = ~n8145 & n16900;
  assign n16902 = ~n9307 & n16901;
  assign n16903 = ~n10554 & n16902;
  assign n16904 = ~n11959 & n16903;
  assign n16905 = ~n13493 & n16904;
  assign n16906 = ~n15167 & n16905;
  assign n16907 = ~n16216 & n16906;
  assign n16908 = ~n16220 & n16907;
  assign n16909 = ~n16466 & n16908;
  assign n16910 = n16476 & n16909;
  assign n16911 = ~n16899 & ~n16910;
  assign n16912 = ~n16465 & ~n16911;
  assign n16913 = ~pi011 & ~n5686;
  assign n16914 = ~n5349 & n16913;
  assign n16915 = ~n5808 & n16914;
  assign n16916 = ~n6056 & n16915;
  assign n16917 = ~n7073 & n16916;
  assign n16918 = ~n8179 & n16917;
  assign n16919 = ~n9344 & n16918;
  assign n16920 = ~n16418 & n16919;
  assign n16921 = ~n16361 & n16920;
  assign n16922 = ~n10594 & n16921;
  assign n16923 = ~n12005 & n16922;
  assign n16924 = ~n13558 & n16923;
  assign n16925 = ~n16216 & n16924;
  assign n16926 = ~n16215 & n16925;
  assign n16927 = n16432 & n16926;
  assign n16928 = n16435 & n16927;
  assign n16929 = n16439 & n16928;
  assign n16930 = n16305 & n16929;
  assign n16931 = n16464 & n16930;
  assign n16932 = ~n15239 & n15275;
  assign n16933 = ~n15061 & n15274;
  assign n16934 = n15266 & ~n16255;
  assign n16935 = ~n16933 & ~n16934;
  assign n16936 = ~n16932 & n16935;
  assign n16937 = n15267 & ~n16285;
  assign n16938 = ~n16216 & n16221;
  assign n16939 = ~n16215 & ~n16220;
  assign n16940 = n16938 & n16939;
  assign n16941 = ~n16937 & n16940;
  assign n16942 = ~n15153 & n15270;
  assign n16943 = ~n14848 & n15265;
  assign n16944 = ~n16942 & ~n16943;
  assign n16945 = n16941 & n16944;
  assign n16946 = n16936 & n16945;
  assign n16947 = ~n16931 & ~n16946;
  assign n16948 = ~n16912 & n16947;
  assign n16949 = n15281 & ~n15419;
  assign n16950 = ~n14741 & n15283;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = n15314 & ~n15616;
  assign n16953 = n15282 & ~n15465;
  assign n16954 = ~n16952 & ~n16953;
  assign n16955 = n16951 & n16954;
  assign n16956 = n6584 & ~n16360;
  assign n16957 = n6643 & ~n16417;
  assign n16958 = ~n6784 & n12054;
  assign n16959 = ~n7158 & n16958;
  assign n16960 = ~n8250 & n16959;
  assign n16961 = ~n9414 & n16960;
  assign n16962 = ~n16957 & n16961;
  assign n16963 = ~n16956 & n16962;
  assign n16964 = ~n10667 & n16963;
  assign n16965 = ~n12083 & n16964;
  assign n16966 = ~n13644 & n16965;
  assign n16967 = ~n16216 & n16966;
  assign n16968 = ~n16215 & n16967;
  assign n16969 = n16222 & n16968;
  assign n16970 = n15301 & ~n15586;
  assign n16971 = ~n15330 & ~n16970;
  assign n16972 = n16969 & n16971;
  assign n16973 = n15287 & ~n15855;
  assign n16974 = n15309 & ~n15886;
  assign n16975 = ~n16973 & ~n16974;
  assign n16976 = n16972 & n16975;
  assign n16977 = n16955 & n16976;
  assign n16978 = n15317 & ~n15657;
  assign n16979 = n15311 & ~n16285;
  assign n16980 = ~n16978 & ~n16979;
  assign n16981 = ~n14848 & n15321;
  assign n16982 = ~n15061 & n15325;
  assign n16983 = ~n16981 & ~n16982;
  assign n16984 = n16980 & n16983;
  assign n16985 = ~n15239 & n15315;
  assign n16986 = ~n14716 & n15286;
  assign n16987 = ~n16985 & ~n16986;
  assign n16988 = n15310 & ~n15536;
  assign n16989 = n15324 & ~n15482;
  assign n16990 = ~n16988 & ~n16989;
  assign n16991 = n16987 & n16990;
  assign n16992 = n15318 & ~n15385;
  assign n16993 = ~n15153 & n15322;
  assign n16994 = ~n16992 & ~n16993;
  assign n16995 = n15304 & ~n15693;
  assign n16996 = n15305 & ~n16255;
  assign n16997 = ~n16995 & ~n16996;
  assign n16998 = n16994 & n16997;
  assign n16999 = n16991 & n16998;
  assign n17000 = n16984 & n16999;
  assign n17001 = n16977 & n17000;
  assign n17002 = ~n15278 & n15331;
  assign n17003 = ~n16216 & n17002;
  assign n17004 = n16939 & n17003;
  assign n17005 = ~n16937 & n17004;
  assign n17006 = n16944 & n17005;
  assign n17007 = n16936 & n17006;
  assign n17008 = ~n17001 & ~n17007;
  assign n17009 = ~n16948 & n17008;
  assign n17010 = n15339 & ~n15465;
  assign n17011 = ~n14741 & n15341;
  assign n17012 = ~n17010 & ~n17011;
  assign n17013 = n15340 & ~n15586;
  assign n17014 = n15359 & ~n15616;
  assign n17015 = ~n17013 & ~n17014;
  assign n17016 = n17012 & n17015;
  assign n17017 = n7475 & ~n16360;
  assign n17018 = n7692 & ~n16417;
  assign n17019 = ~n7505 & ~n7663;
  assign n17020 = ~n7869 & n17019;
  assign n17021 = ~n8346 & n17020;
  assign n17022 = ~n9485 & n17021;
  assign n17023 = ~n17018 & n17022;
  assign n17024 = ~n17017 & n17023;
  assign n17025 = ~n10741 & n17024;
  assign n17026 = ~n12158 & n17025;
  assign n17027 = ~n13693 & n17026;
  assign n17028 = ~n16216 & n17027;
  assign n17029 = ~n16215 & n17028;
  assign n17030 = n16222 & n17029;
  assign n17031 = ~n15385 & ~n16209;
  assign n17032 = n17030 & n17031;
  assign n17033 = n15364 & ~n15886;
  assign n17034 = n15345 & ~n15855;
  assign n17035 = ~n17033 & ~n17034;
  assign n17036 = n17032 & n17035;
  assign n17037 = n17016 & n17036;
  assign n17038 = ~n15330 & n15369;
  assign n17039 = ~n14848 & n15373;
  assign n17040 = ~n17038 & ~n17039;
  assign n17041 = ~n15061 & n15365;
  assign n17042 = n15370 & ~n15482;
  assign n17043 = ~n17041 & ~n17042;
  assign n17044 = n17040 & n17043;
  assign n17045 = ~n14716 & n15344;
  assign n17046 = ~n15239 & n15380;
  assign n17047 = ~n17045 & ~n17046;
  assign n17048 = n15372 & ~n15657;
  assign n17049 = ~n15153 & n15360;
  assign n17050 = ~n17048 & ~n17049;
  assign n17051 = n17047 & n17050;
  assign n17052 = n15376 & ~n16255;
  assign n17053 = n15377 & ~n15693;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = n15366 & ~n16285;
  assign n17056 = n15379 & ~n15536;
  assign n17057 = ~n17055 & ~n17056;
  assign n17058 = n17054 & n17057;
  assign n17059 = n17051 & n17058;
  assign n17060 = n17044 & n17059;
  assign n17061 = n17037 & n17060;
  assign n17062 = ~n6401 & n10675;
  assign n17063 = ~n6784 & n17062;
  assign n17064 = ~n7158 & n17063;
  assign n17065 = ~n8250 & n17064;
  assign n17066 = ~n9414 & n17065;
  assign n17067 = ~n16957 & n17066;
  assign n17068 = ~n16956 & n17067;
  assign n17069 = ~n10667 & n17068;
  assign n17070 = ~n12083 & n17069;
  assign n17071 = ~n13644 & n17070;
  assign n17072 = ~n16216 & n17071;
  assign n17073 = ~n16215 & n17072;
  assign n17074 = n16222 & n17073;
  assign n17075 = n16971 & n17074;
  assign n17076 = n16975 & n17075;
  assign n17077 = n16955 & n17076;
  assign n17078 = n17000 & n17077;
  assign n17079 = n15415 & ~n16255;
  assign n17080 = ~n14848 & n15412;
  assign n17081 = ~n15061 & n15403;
  assign n17082 = ~n17080 & ~n17081;
  assign n17083 = ~n17079 & n17082;
  assign n17084 = n14455 & ~n16216;
  assign n17085 = ~n15419 & n17084;
  assign n17086 = ~n16221 & n16939;
  assign n17087 = n17085 & n17086;
  assign n17088 = ~n15239 & n15404;
  assign n17089 = ~n15153 & n15405;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = ~n15330 & n15414;
  assign n17092 = n15411 & ~n16285;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = n17090 & n17093;
  assign n17095 = n17087 & n17094;
  assign n17096 = n17083 & n17095;
  assign n17097 = ~n17078 & ~n17096;
  assign n17098 = ~n17061 & n17097;
  assign n17099 = ~n17009 & n17098;
  assign n17100 = ~n7505 & n8357;
  assign n17101 = ~n7869 & n17100;
  assign n17102 = ~n8346 & n17101;
  assign n17103 = ~n9485 & n17102;
  assign n17104 = ~n17018 & n17103;
  assign n17105 = ~n17017 & n17104;
  assign n17106 = ~n10741 & n17105;
  assign n17107 = ~n12158 & n17106;
  assign n17108 = ~n13693 & n17107;
  assign n17109 = ~n16216 & n17108;
  assign n17110 = ~n16215 & n17109;
  assign n17111 = n16222 & n17110;
  assign n17112 = n17031 & n17111;
  assign n17113 = n17035 & n17112;
  assign n17114 = n17016 & n17113;
  assign n17115 = n17060 & n17114;
  assign n17116 = n15461 & ~n16255;
  assign n17117 = ~n15153 & n15458;
  assign n17118 = ~n17116 & ~n17117;
  assign n17119 = ~n14848 & n15457;
  assign n17120 = ~n15061 & n15450;
  assign n17121 = ~n17119 & ~n17120;
  assign n17122 = n17118 & n17121;
  assign n17123 = n14454 & ~n16216;
  assign n17124 = ~n15465 & n17123;
  assign n17125 = ~n16209 & n17124;
  assign n17126 = n17086 & n17125;
  assign n17127 = ~n15239 & n15460;
  assign n17128 = n15447 & ~n16285;
  assign n17129 = ~n17127 & ~n17128;
  assign n17130 = ~n15330 & n15449;
  assign n17131 = ~n15385 & n15446;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = n17129 & n17132;
  assign n17134 = n17126 & n17133;
  assign n17135 = n17122 & n17134;
  assign n17136 = ~n13726 & n15440;
  assign n17137 = ~n16216 & n17136;
  assign n17138 = ~n15419 & n17137;
  assign n17139 = n17086 & n17138;
  assign n17140 = n17094 & n17139;
  assign n17141 = n17083 & n17140;
  assign n17142 = ~n17135 & ~n17141;
  assign n17143 = ~n17115 & n17142;
  assign n17144 = ~n17099 & n17143;
  assign n17145 = n14743 & ~n15586;
  assign n17146 = ~n16211 & ~n17145;
  assign n17147 = ~n14741 & n14742;
  assign n17148 = n14762 & ~n15616;
  assign n17149 = ~n17147 & ~n17148;
  assign n17150 = n17146 & n17149;
  assign n17151 = n8574 & ~n16360;
  assign n17152 = n8484 & ~n16417;
  assign n17153 = ~n8834 & n11377;
  assign n17154 = ~n10002 & n17153;
  assign n17155 = ~n17152 & n17154;
  assign n17156 = ~n17151 & n17155;
  assign n17157 = ~n11297 & n17156;
  assign n17158 = ~n12240 & n17157;
  assign n17159 = ~n13135 & n17158;
  assign n17160 = ~n16216 & n17159;
  assign n17161 = ~n16215 & n17160;
  assign n17162 = n16222 & n17161;
  assign n17163 = ~n15482 & ~n16209;
  assign n17164 = n17162 & n17163;
  assign n17165 = n14767 & ~n15886;
  assign n17166 = n14747 & ~n15855;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = n17164 & n17167;
  assign n17169 = n17150 & n17168;
  assign n17170 = n14782 & ~n15536;
  assign n17171 = n14776 & ~n14848;
  assign n17172 = ~n17170 & ~n17171;
  assign n17173 = n14769 & ~n16285;
  assign n17174 = n14763 & ~n15153;
  assign n17175 = ~n17173 & ~n17174;
  assign n17176 = n17172 & n17175;
  assign n17177 = n14783 & ~n15239;
  assign n17178 = ~n14716 & n14746;
  assign n17179 = ~n17177 & ~n17178;
  assign n17180 = n14768 & ~n15061;
  assign n17181 = n14773 & ~n15330;
  assign n17182 = ~n17180 & ~n17181;
  assign n17183 = n17179 & n17182;
  assign n17184 = n14780 & ~n15693;
  assign n17185 = n14772 & ~n15385;
  assign n17186 = ~n17184 & ~n17185;
  assign n17187 = n14775 & ~n15657;
  assign n17188 = n14779 & ~n16255;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = n17186 & n17189;
  assign n17191 = n17183 & n17190;
  assign n17192 = n17176 & n17191;
  assign n17193 = n17169 & n17192;
  assign n17194 = ~n13764 & n15483;
  assign n17195 = ~n16216 & n17194;
  assign n17196 = ~n15465 & n17195;
  assign n17197 = ~n16209 & n17196;
  assign n17198 = n17086 & n17197;
  assign n17199 = n17133 & n17198;
  assign n17200 = n17122 & n17199;
  assign n17201 = ~n17193 & ~n17200;
  assign n17202 = ~n17144 & n17201;
  assign n17203 = pi017 & ~n8633;
  assign n17204 = ~n8455 & n17203;
  assign n17205 = ~n8834 & n17204;
  assign n17206 = ~n10002 & n17205;
  assign n17207 = ~n17152 & n17206;
  assign n17208 = ~n17151 & n17207;
  assign n17209 = ~n11297 & n17208;
  assign n17210 = ~n12240 & n17209;
  assign n17211 = ~n13135 & n17210;
  assign n17212 = ~n16216 & n17211;
  assign n17213 = ~n16215 & n17212;
  assign n17214 = n16222 & n17213;
  assign n17215 = n17163 & n17214;
  assign n17216 = n17167 & n17215;
  assign n17217 = n17150 & n17216;
  assign n17218 = n17192 & n17217;
  assign n17219 = n14735 & ~n15153;
  assign n17220 = n14724 & ~n14848;
  assign n17221 = ~n17219 & ~n17220;
  assign n17222 = n14717 & ~n15061;
  assign n17223 = n14720 & ~n15239;
  assign n17224 = ~n17222 & ~n17223;
  assign n17225 = n17221 & n17224;
  assign n17226 = n14728 & ~n16255;
  assign n17227 = n14721 & ~n15330;
  assign n17228 = ~n17226 & ~n17227;
  assign n17229 = n14727 & ~n16285;
  assign n17230 = n14725 & ~n15385;
  assign n17231 = ~n17229 & ~n17230;
  assign n17232 = n17228 & n17231;
  assign n17233 = n14452 & ~n16216;
  assign n17234 = ~n14741 & n17233;
  assign n17235 = ~n16209 & n17234;
  assign n17236 = ~n16211 & n17235;
  assign n17237 = n14718 & ~n15482;
  assign n17238 = n17086 & ~n17237;
  assign n17239 = n17236 & n17238;
  assign n17240 = n17232 & n17239;
  assign n17241 = n17225 & n17240;
  assign n17242 = ~n17218 & ~n17241;
  assign n17243 = ~n17202 & n17242;
  assign n17244 = ~pi018 & ~n8900;
  assign n17245 = ~n9533 & n17244;
  assign n17246 = ~n10787 & n17245;
  assign n17247 = ~n11611 & n17246;
  assign n17248 = ~n13820 & n17247;
  assign n17249 = ~n16216 & n17248;
  assign n17250 = ~n14741 & n17249;
  assign n17251 = ~n16209 & n17250;
  assign n17252 = ~n16211 & n17251;
  assign n17253 = n17238 & n17252;
  assign n17254 = n17232 & n17253;
  assign n17255 = n17225 & n17254;
  assign n17256 = ~n17243 & ~n17255;
  assign n17257 = ~n16209 & ~n16211;
  assign n17258 = n15494 & ~n15586;
  assign n17259 = n15531 & ~n15616;
  assign n17260 = ~n17258 & ~n17259;
  assign n17261 = n17257 & n17260;
  assign n17262 = n9793 & ~n16360;
  assign n17263 = n9854 & ~n16417;
  assign n17264 = ~n9929 & n11562;
  assign n17265 = ~n17263 & n17264;
  assign n17266 = ~n17262 & n17265;
  assign n17267 = ~n11266 & n17266;
  assign n17268 = ~n11588 & n17267;
  assign n17269 = ~n13859 & n17268;
  assign n17270 = ~n16216 & n17269;
  assign n17271 = ~n16215 & n17270;
  assign n17272 = n16222 & n17271;
  assign n17273 = ~n15536 & ~n16208;
  assign n17274 = n17272 & n17273;
  assign n17275 = ~n15239 & n15516;
  assign n17276 = ~n14716 & n15496;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = n17274 & n17277;
  assign n17279 = n17261 & n17278;
  assign n17280 = n15510 & ~n15693;
  assign n17281 = ~n15385 & n15511;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = ~n15061 & n15530;
  assign n17284 = ~n15482 & n15520;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = n17282 & n17285;
  assign n17287 = ~n15153 & n15523;
  assign n17288 = n15524 & ~n15657;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = ~n15330 & n15528;
  assign n17291 = n15517 & ~n16285;
  assign n17292 = ~n17290 & ~n17291;
  assign n17293 = n17289 & n17292;
  assign n17294 = n15497 & ~n15855;
  assign n17295 = n15515 & ~n15886;
  assign n17296 = ~n17294 & ~n17295;
  assign n17297 = n15527 & ~n16255;
  assign n17298 = ~n14848 & n15521;
  assign n17299 = ~n17297 & ~n17298;
  assign n17300 = n17296 & n17299;
  assign n17301 = n17293 & n17300;
  assign n17302 = n17286 & n17301;
  assign n17303 = n17279 & n17302;
  assign n17304 = ~n17256 & ~n17303;
  assign n17305 = ~n9763 & n15547;
  assign n17306 = ~n9929 & n17305;
  assign n17307 = ~n17263 & n17306;
  assign n17308 = ~n17262 & n17307;
  assign n17309 = ~n11266 & n17308;
  assign n17310 = ~n11588 & n17309;
  assign n17311 = ~n13859 & n17310;
  assign n17312 = ~n16216 & n17311;
  assign n17313 = ~n16215 & n17312;
  assign n17314 = n16222 & n17313;
  assign n17315 = n17273 & n17314;
  assign n17316 = n17277 & n17315;
  assign n17317 = n17261 & n17316;
  assign n17318 = n17302 & n17317;
  assign n17319 = n14451 & ~n16216;
  assign n17320 = ~n15586 & n17319;
  assign n17321 = ~n16208 & n17320;
  assign n17322 = n17257 & n17321;
  assign n17323 = ~n15482 & n15575;
  assign n17324 = n17086 & ~n17323;
  assign n17325 = ~n15536 & n15578;
  assign n17326 = n15574 & ~n16255;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = n17324 & n17327;
  assign n17329 = n17322 & n17328;
  assign n17330 = ~n15385 & n15568;
  assign n17331 = ~n14848 & n15573;
  assign n17332 = ~n15239 & n15579;
  assign n17333 = ~n17331 & ~n17332;
  assign n17334 = ~n17330 & n17333;
  assign n17335 = n15581 & ~n16285;
  assign n17336 = ~n15153 & n15566;
  assign n17337 = ~n17335 & ~n17336;
  assign n17338 = ~n15061 & n15582;
  assign n17339 = ~n15330 & n15569;
  assign n17340 = ~n17338 & ~n17339;
  assign n17341 = n17337 & n17340;
  assign n17342 = n17334 & n17341;
  assign n17343 = n17329 & n17342;
  assign n17344 = ~n15061 & n15588;
  assign n17345 = n15603 & ~n16255;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = n15605 & ~n16285;
  assign n17348 = ~n15536 & n15604;
  assign n17349 = ~n17347 & ~n17348;
  assign n17350 = n17346 & n17349;
  assign n17351 = n16210 & ~n16211;
  assign n17352 = n14577 & ~n16216;
  assign n17353 = ~n15616 & n17352;
  assign n17354 = ~n16224 & n17353;
  assign n17355 = n17086 & n17354;
  assign n17356 = n17351 & n17355;
  assign n17357 = n17350 & n17356;
  assign n17358 = ~n14848 & n15608;
  assign n17359 = ~n15239 & n15609;
  assign n17360 = ~n15385 & n15587;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = ~n17358 & n17361;
  assign n17363 = ~n15482 & n15611;
  assign n17364 = ~n15330 & n15590;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = n15612 & ~n15657;
  assign n17367 = ~n15153 & n15591;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = n17365 & n17368;
  assign n17370 = n17362 & n17369;
  assign n17371 = n17357 & n17370;
  assign n17372 = ~n17343 & ~n17371;
  assign n17373 = ~n17318 & n17372;
  assign n17374 = ~n15616 & n15649;
  assign n17375 = ~n16211 & ~n17374;
  assign n17376 = n16210 & n17375;
  assign n17377 = n11103 & ~n16360;
  assign n17378 = n11072 & ~n16417;
  assign n17379 = ~n11188 & n12317;
  assign n17380 = ~n17378 & n17379;
  assign n17381 = ~n17377 & n17380;
  assign n17382 = ~n12380 & n17381;
  assign n17383 = ~n14045 & n17382;
  assign n17384 = ~n16216 & n17383;
  assign n17385 = ~n16215 & n17384;
  assign n17386 = n16222 & n17385;
  assign n17387 = ~n15657 & ~n16224;
  assign n17388 = n17386 & n17387;
  assign n17389 = n15620 & ~n15855;
  assign n17390 = n15651 & ~n15886;
  assign n17391 = ~n17389 & ~n17390;
  assign n17392 = n17388 & n17391;
  assign n17393 = n17376 & n17392;
  assign n17394 = n15641 & ~n16285;
  assign n17395 = ~n15239 & n15645;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = ~n15536 & n15648;
  assign n17398 = ~n15385 & n15638;
  assign n17399 = ~n17397 & ~n17398;
  assign n17400 = n17396 & n17399;
  assign n17401 = ~n15482 & n15636;
  assign n17402 = ~n14716 & n15619;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~n15330 & n15652;
  assign n17405 = n15644 & ~n15693;
  assign n17406 = ~n17404 & ~n17405;
  assign n17407 = n17403 & n17406;
  assign n17408 = n15632 & ~n16255;
  assign n17409 = ~n14848 & n15637;
  assign n17410 = ~n17408 & ~n17409;
  assign n17411 = ~n15061 & n15631;
  assign n17412 = ~n15153 & n15642;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = n17410 & n17413;
  assign n17415 = n17407 & n17414;
  assign n17416 = n17400 & n17415;
  assign n17417 = n17393 & n17416;
  assign n17418 = n12841 & ~n16360;
  assign n17419 = n12713 & ~n16417;
  assign n17420 = n12774 & ~n12902;
  assign n17421 = ~n17419 & n17420;
  assign n17422 = ~n17418 & n17421;
  assign n17423 = ~n14009 & n17422;
  assign n17424 = ~n16216 & n17423;
  assign n17425 = ~n16215 & n17424;
  assign n17426 = n16222 & n17425;
  assign n17427 = ~n15693 & ~n16224;
  assign n17428 = n17426 & n17427;
  assign n17429 = ~n15061 & n15685;
  assign n17430 = ~n15153 & n15684;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = n17428 & n17431;
  assign n17433 = n16214 & n17432;
  assign n17434 = n15674 & ~n15886;
  assign n17435 = ~n14716 & n15659;
  assign n17436 = ~n17434 & ~n17435;
  assign n17437 = ~n15385 & n15677;
  assign n17438 = ~n15536 & n15678;
  assign n17439 = ~n17437 & ~n17438;
  assign n17440 = n17436 & n17439;
  assign n17441 = n15688 & ~n16255;
  assign n17442 = ~n15330 & n15672;
  assign n17443 = ~n17441 & ~n17442;
  assign n17444 = n15680 & ~n16285;
  assign n17445 = ~n14848 & n15681;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = n17443 & n17446;
  assign n17448 = ~n15239 & n15668;
  assign n17449 = ~n15482 & n15673;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = n15658 & ~n15855;
  assign n17452 = ~n15657 & n15687;
  assign n17453 = ~n17451 & ~n17452;
  assign n17454 = n17450 & n17453;
  assign n17455 = n17447 & n17454;
  assign n17456 = n17440 & n17455;
  assign n17457 = n17433 & n17456;
  assign n17458 = ~n17417 & ~n17457;
  assign n17459 = n17373 & n17458;
  assign n17460 = ~n17304 & n17459;
  assign n17461 = ~n11042 & n15697;
  assign n17462 = ~n11188 & n17461;
  assign n17463 = ~n17378 & n17462;
  assign n17464 = ~n17377 & n17463;
  assign n17465 = ~n12380 & n17464;
  assign n17466 = ~n14045 & n17465;
  assign n17467 = ~n16216 & n17466;
  assign n17468 = ~n16215 & n17467;
  assign n17469 = n16222 & n17468;
  assign n17470 = n17387 & n17469;
  assign n17471 = n17391 & n17470;
  assign n17472 = n17376 & n17471;
  assign n17473 = n17416 & n17472;
  assign n17474 = pi023 & ~n12743;
  assign n17475 = ~n12773 & n17474;
  assign n17476 = ~n12902 & n17475;
  assign n17477 = ~n17419 & n17476;
  assign n17478 = ~n17418 & n17477;
  assign n17479 = ~n14009 & n17478;
  assign n17480 = ~n16216 & n17479;
  assign n17481 = ~n16215 & n17480;
  assign n17482 = n16222 & n17481;
  assign n17483 = n17427 & n17482;
  assign n17484 = n17431 & n17483;
  assign n17485 = n16214 & n17484;
  assign n17486 = n17456 & n17485;
  assign n17487 = ~n13906 & n15723;
  assign n17488 = ~n16216 & n17487;
  assign n17489 = ~n15586 & n17488;
  assign n17490 = ~n16208 & n17489;
  assign n17491 = n17257 & n17490;
  assign n17492 = n17328 & n17491;
  assign n17493 = n17342 & n17492;
  assign n17494 = ~n14073 & n15730;
  assign n17495 = ~n16216 & n17494;
  assign n17496 = ~n15616 & n17495;
  assign n17497 = ~n16224 & n17496;
  assign n17498 = n17086 & n17497;
  assign n17499 = n17351 & n17498;
  assign n17500 = n17350 & n17499;
  assign n17501 = n17370 & n17500;
  assign n17502 = ~n17493 & ~n17501;
  assign n17503 = ~n17486 & n17502;
  assign n17504 = ~n17473 & n17503;
  assign n17505 = ~n17460 & n17504;
  assign n17506 = ~n15385 & n15881;
  assign n17507 = ~n15657 & n15867;
  assign n17508 = ~n17506 & ~n17507;
  assign n17509 = ~n15693 & n15861;
  assign n17510 = ~n14848 & n15873;
  assign n17511 = ~n17509 & ~n17510;
  assign n17512 = n17508 & n17511;
  assign n17513 = n14676 & ~n16216;
  assign n17514 = ~n16215 & n17513;
  assign n17515 = n16222 & n17514;
  assign n17516 = ~n15886 & ~n16224;
  assign n17517 = n17515 & n17516;
  assign n17518 = n16214 & n17517;
  assign n17519 = n17512 & n17518;
  assign n17520 = n15874 & ~n16285;
  assign n17521 = n15870 & ~n16255;
  assign n17522 = ~n17520 & ~n17521;
  assign n17523 = ~n15153 & n15877;
  assign n17524 = ~n15239 & n15878;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = n17522 & n17525;
  assign n17527 = ~n15482 & n15871;
  assign n17528 = ~n15330 & n15866;
  assign n17529 = ~n17527 & ~n17528;
  assign n17530 = ~n15061 & n15865;
  assign n17531 = ~n15536 & n15880;
  assign n17532 = ~n17530 & ~n17531;
  assign n17533 = n17529 & n17532;
  assign n17534 = n17526 & n17533;
  assign n17535 = n17519 & n17534;
  assign n17536 = n14416 & ~n16417;
  assign n17537 = n14320 & ~n16360;
  assign n17538 = ~n14519 & n15744;
  assign n17539 = ~n17537 & n17538;
  assign n17540 = ~n17536 & n17539;
  assign n17541 = ~n16216 & n17540;
  assign n17542 = ~n16215 & n17541;
  assign n17543 = n16222 & n17542;
  assign n17544 = ~n15855 & ~n16224;
  assign n17545 = n17543 & n17544;
  assign n17546 = ~n14848 & n15845;
  assign n17547 = ~n16232 & ~n17546;
  assign n17548 = n17545 & n17547;
  assign n17549 = n16214 & n17548;
  assign n17550 = ~n15657 & n15781;
  assign n17551 = n15823 & ~n16255;
  assign n17552 = ~n17550 & ~n17551;
  assign n17553 = ~n15239 & n15791;
  assign n17554 = ~n15061 & n15811;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 = n17552 & n17555;
  assign n17557 = ~n14716 & n15742;
  assign n17558 = ~n15330 & n15778;
  assign n17559 = ~n17557 & ~n17558;
  assign n17560 = ~n15385 & n15833;
  assign n17561 = ~n15153 & n15800;
  assign n17562 = ~n17560 & ~n17561;
  assign n17563 = n17559 & n17562;
  assign n17564 = n15771 & ~n16285;
  assign n17565 = ~n15536 & n15755;
  assign n17566 = ~n17564 & ~n17565;
  assign n17567 = ~n15693 & n15827;
  assign n17568 = ~n15482 & n15850;
  assign n17569 = ~n17567 & ~n17568;
  assign n17570 = n17566 & n17569;
  assign n17571 = n17563 & n17570;
  assign n17572 = n17556 & n17571;
  assign n17573 = n17549 & n17572;
  assign n17574 = ~n17535 & ~n17573;
  assign n17575 = ~n17505 & n17574;
  assign n17576 = ~n14568 & ~n16216;
  assign n17577 = ~n16215 & n17576;
  assign n17578 = n16222 & n17577;
  assign n17579 = n16225 & n17578;
  assign n17580 = n16229 & n17579;
  assign n17581 = n16214 & n17580;
  assign n17582 = n16297 & n17581;
  assign n17583 = pi025 & ~n14350;
  assign n17584 = ~n14381 & n17583;
  assign n17585 = ~n14519 & n17584;
  assign n17586 = ~n17537 & n17585;
  assign n17587 = ~n17536 & n17586;
  assign n17588 = ~n16216 & n17587;
  assign n17589 = ~n16215 & n17588;
  assign n17590 = n16222 & n17589;
  assign n17591 = n17544 & n17590;
  assign n17592 = n17547 & n17591;
  assign n17593 = n16214 & n17592;
  assign n17594 = n17572 & n17593;
  assign n17595 = ~n13093 & n14118;
  assign n17596 = ~n16216 & n17595;
  assign n17597 = ~n16215 & n17596;
  assign n17598 = n16222 & n17597;
  assign n17599 = n17516 & n17598;
  assign n17600 = n16214 & n17599;
  assign n17601 = n17512 & n17600;
  assign n17602 = n17534 & n17601;
  assign n17603 = ~n17594 & ~n17602;
  assign n17604 = ~n17582 & n17603;
  assign n17605 = ~n17575 & n17604;
  assign n17606 = ~n16298 & ~n17605;
  assign n17607 = ~n2572 & ~n3066;
  assign n17608 = ~n3983 & n17607;
  assign n17609 = ~n4024 & n17608;
  assign n17610 = ~n4999 & n17609;
  assign n17611 = ~n5827 & n17610;
  assign n17612 = ~n6893 & n17611;
  assign n17613 = ~n7890 & n17612;
  assign n17614 = ~n9131 & n17613;
  assign n17615 = ~n10278 & n17614;
  assign n17616 = ~n11662 & n17615;
  assign n17617 = ~n13191 & n17616;
  assign n17618 = ~n14848 & n17617;
  assign n17619 = ~n16232 & ~n17618;
  assign n17620 = ~n12841 & ~n12902;
  assign n17621 = ~n14009 & n17620;
  assign n17622 = ~n15693 & n17621;
  assign n17623 = ~n11103 & ~n11188;
  assign n17624 = ~n12380 & n17623;
  assign n17625 = ~n14045 & n17624;
  assign n17626 = ~n15657 & n17625;
  assign n17627 = ~n17622 & ~n17626;
  assign n17628 = n17619 & n17627;
  assign n17629 = ~n16212 & n17257;
  assign n17630 = n16176 & ~n16417;
  assign n17631 = ~n16144 & ~n16175;
  assign n17632 = ~n16360 & n17631;
  assign n17633 = ~n17630 & n17632;
  assign n17634 = ~n16216 & n17633;
  assign n17635 = ~n16215 & n17634;
  assign n17636 = n16222 & n17635;
  assign n17637 = ~n16208 & ~n16224;
  assign n17638 = n17636 & n17637;
  assign n17639 = n17629 & n17638;
  assign n17640 = n17628 & n17639;
  assign n17641 = ~n14320 & ~n14519;
  assign n17642 = ~n15855 & n17641;
  assign n17643 = ~n14568 & ~n14716;
  assign n17644 = ~n8574 & ~n8834;
  assign n17645 = ~n10002 & n17644;
  assign n17646 = ~n11297 & n17645;
  assign n17647 = ~n12240 & n17646;
  assign n17648 = ~n13135 & n17647;
  assign n17649 = ~n15482 & n17648;
  assign n17650 = ~n17643 & ~n17649;
  assign n17651 = ~n17642 & n17650;
  assign n17652 = ~n1587 & ~n2242;
  assign n17653 = ~n3095 & n17652;
  assign n17654 = ~n3997 & n17653;
  assign n17655 = ~n4837 & n17654;
  assign n17656 = ~n5822 & n17655;
  assign n17657 = ~n6820 & n17656;
  assign n17658 = ~n7785 & n17657;
  assign n17659 = ~n9027 & n17658;
  assign n17660 = ~n10245 & n17659;
  assign n17661 = ~n11536 & n17660;
  assign n17662 = ~n13036 & n17661;
  assign n17663 = ~n14653 & n17662;
  assign n17664 = ~n16255 & n17663;
  assign n17665 = ~n7475 & ~n7869;
  assign n17666 = ~n8346 & n17665;
  assign n17667 = ~n9485 & n17666;
  assign n17668 = ~n10741 & n17667;
  assign n17669 = ~n12158 & n17668;
  assign n17670 = ~n13693 & n17669;
  assign n17671 = ~n15385 & n17670;
  assign n17672 = ~n17664 & ~n17671;
  assign n17673 = ~n6584 & ~n6784;
  assign n17674 = ~n7158 & n17673;
  assign n17675 = ~n8250 & n17674;
  assign n17676 = ~n9414 & n17675;
  assign n17677 = ~n10667 & n17676;
  assign n17678 = ~n12083 & n17677;
  assign n17679 = ~n13644 & n17678;
  assign n17680 = ~n15330 & n17679;
  assign n17681 = ~n3620 & ~n3940;
  assign n17682 = ~n4001 & n17681;
  assign n17683 = ~n5043 & n17682;
  assign n17684 = ~n5943 & n17683;
  assign n17685 = ~n6951 & n17684;
  assign n17686 = ~n8037 & n17685;
  assign n17687 = ~n9200 & n17686;
  assign n17688 = ~n10445 & n17687;
  assign n17689 = ~n11846 & n17688;
  assign n17690 = ~n13393 & n17689;
  assign n17691 = ~n15061 & n17690;
  assign n17692 = ~n17680 & ~n17691;
  assign n17693 = n17672 & n17692;
  assign n17694 = ~n9793 & ~n9929;
  assign n17695 = ~n11266 & n17694;
  assign n17696 = ~n11588 & n17695;
  assign n17697 = ~n13859 & n17696;
  assign n17698 = ~n15536 & n17697;
  assign n17699 = ~n5657 & ~n5808;
  assign n17700 = ~n6056 & n17699;
  assign n17701 = ~n7073 & n17700;
  assign n17702 = ~n8179 & n17701;
  assign n17703 = ~n9344 & n17702;
  assign n17704 = ~n10594 & n17703;
  assign n17705 = ~n12005 & n17704;
  assign n17706 = ~n13558 & n17705;
  assign n17707 = ~n15239 & n17706;
  assign n17708 = ~n17698 & ~n17707;
  assign n17709 = ~n750 & ~n1372;
  assign n17710 = ~n2243 & n17709;
  assign n17711 = ~n3104 & n17710;
  assign n17712 = ~n3971 & n17711;
  assign n17713 = ~n4872 & n17712;
  assign n17714 = ~n5801 & n17713;
  assign n17715 = ~n6739 & n17714;
  assign n17716 = ~n7807 & n17715;
  assign n17717 = ~n8989 & n17716;
  assign n17718 = ~n10273 & n17717;
  assign n17719 = ~n11499 & n17718;
  assign n17720 = ~n13076 & n17719;
  assign n17721 = ~n14698 & n17720;
  assign n17722 = ~n16285 & n17721;
  assign n17723 = ~n4489 & ~n4817;
  assign n17724 = ~n4902 & n17723;
  assign n17725 = ~n6001 & n17724;
  assign n17726 = ~n7014 & n17725;
  assign n17727 = ~n8114 & n17726;
  assign n17728 = ~n9276 & n17727;
  assign n17729 = ~n10523 & n17728;
  assign n17730 = ~n11928 & n17729;
  assign n17731 = ~n13479 & n17730;
  assign n17732 = ~n15153 & n17731;
  assign n17733 = ~n17722 & ~n17732;
  assign n17734 = n17708 & n17733;
  assign n17735 = n17693 & n17734;
  assign n17736 = n17651 & n17735;
  assign n17737 = n17640 & n17736;
  assign n17738 = ~n17606 & ~n17737;
  assign n17739 = ~pi027 & ~n16144;
  assign n17740 = ~n16175 & n17739;
  assign n17741 = ~n16360 & n17740;
  assign n17742 = ~n17630 & n17741;
  assign n17743 = ~n16216 & n17742;
  assign n17744 = ~n16215 & n17743;
  assign n17745 = n16222 & n17744;
  assign n17746 = n17637 & n17745;
  assign n17747 = n17629 & n17746;
  assign n17748 = n17628 & n17747;
  assign n17749 = n17736 & n17748;
  assign n17750 = ~n16232 & ~n17643;
  assign n17751 = ~n9854 & ~n9929;
  assign n17752 = ~n11266 & n17751;
  assign n17753 = ~n11588 & n17752;
  assign n17754 = ~n13859 & n17753;
  assign n17755 = ~n15536 & n17754;
  assign n17756 = ~n6643 & ~n6784;
  assign n17757 = ~n7158 & n17756;
  assign n17758 = ~n8250 & n17757;
  assign n17759 = ~n9414 & n17758;
  assign n17760 = ~n10667 & n17759;
  assign n17761 = ~n12083 & n17760;
  assign n17762 = ~n13644 & n17761;
  assign n17763 = ~n15330 & n17762;
  assign n17764 = ~n17755 & ~n17763;
  assign n17765 = n17750 & n17764;
  assign n17766 = ~n16176 & ~n16360;
  assign n17767 = ~n16417 & ~n17766;
  assign n17768 = ~n16216 & n17767;
  assign n17769 = ~n16215 & n17768;
  assign n17770 = n16222 & n17769;
  assign n17771 = n17637 & n17770;
  assign n17772 = n17629 & n17771;
  assign n17773 = n17765 & n17772;
  assign n17774 = ~n7692 & ~n7869;
  assign n17775 = ~n8346 & n17774;
  assign n17776 = ~n9485 & n17775;
  assign n17777 = ~n10741 & n17776;
  assign n17778 = ~n12158 & n17777;
  assign n17779 = ~n13693 & n17778;
  assign n17780 = ~n15385 & n17779;
  assign n17781 = ~n3591 & ~n3940;
  assign n17782 = ~n4001 & n17781;
  assign n17783 = ~n5043 & n17782;
  assign n17784 = ~n5943 & n17783;
  assign n17785 = ~n6951 & n17784;
  assign n17786 = ~n8037 & n17785;
  assign n17787 = ~n9200 & n17786;
  assign n17788 = ~n10445 & n17787;
  assign n17789 = ~n11846 & n17788;
  assign n17790 = ~n13393 & n17789;
  assign n17791 = ~n15061 & n17790;
  assign n17792 = ~n1740 & ~n2242;
  assign n17793 = ~n3095 & n17792;
  assign n17794 = ~n3997 & n17793;
  assign n17795 = ~n4837 & n17794;
  assign n17796 = ~n5822 & n17795;
  assign n17797 = ~n6820 & n17796;
  assign n17798 = ~n7785 & n17797;
  assign n17799 = ~n9027 & n17798;
  assign n17800 = ~n10245 & n17799;
  assign n17801 = ~n11536 & n17800;
  assign n17802 = ~n13036 & n17801;
  assign n17803 = ~n14653 & n17802;
  assign n17804 = ~n16255 & n17803;
  assign n17805 = ~n17791 & ~n17804;
  assign n17806 = ~n17780 & n17805;
  assign n17807 = ~n12713 & ~n12902;
  assign n17808 = ~n14009 & n17807;
  assign n17809 = ~n15693 & n17808;
  assign n17810 = ~n4430 & ~n4817;
  assign n17811 = ~n4902 & n17810;
  assign n17812 = ~n6001 & n17811;
  assign n17813 = ~n7014 & n17812;
  assign n17814 = ~n8114 & n17813;
  assign n17815 = ~n9276 & n17814;
  assign n17816 = ~n10523 & n17815;
  assign n17817 = ~n11928 & n17816;
  assign n17818 = ~n13479 & n17817;
  assign n17819 = ~n15153 & n17818;
  assign n17820 = ~n17809 & ~n17819;
  assign n17821 = ~n1238 & ~n1372;
  assign n17822 = ~n2243 & n17821;
  assign n17823 = ~n3104 & n17822;
  assign n17824 = ~n3971 & n17823;
  assign n17825 = ~n4872 & n17824;
  assign n17826 = ~n5801 & n17825;
  assign n17827 = ~n6739 & n17826;
  assign n17828 = ~n7807 & n17827;
  assign n17829 = ~n8989 & n17828;
  assign n17830 = ~n10273 & n17829;
  assign n17831 = ~n11499 & n17830;
  assign n17832 = ~n13076 & n17831;
  assign n17833 = ~n14698 & n17832;
  assign n17834 = ~n16285 & n17833;
  assign n17835 = ~n14416 & ~n14519;
  assign n17836 = ~n15855 & n17835;
  assign n17837 = ~n17834 & ~n17836;
  assign n17838 = n17820 & n17837;
  assign n17839 = ~n8484 & ~n8834;
  assign n17840 = ~n10002 & n17839;
  assign n17841 = ~n11297 & n17840;
  assign n17842 = ~n12240 & n17841;
  assign n17843 = ~n13135 & n17842;
  assign n17844 = ~n15482 & n17843;
  assign n17845 = ~n5627 & ~n5808;
  assign n17846 = ~n6056 & n17845;
  assign n17847 = ~n7073 & n17846;
  assign n17848 = ~n8179 & n17847;
  assign n17849 = ~n9344 & n17848;
  assign n17850 = ~n10594 & n17849;
  assign n17851 = ~n12005 & n17850;
  assign n17852 = ~n13558 & n17851;
  assign n17853 = ~n15239 & n17852;
  assign n17854 = ~n17844 & ~n17853;
  assign n17855 = ~n11072 & ~n11188;
  assign n17856 = ~n12380 & n17855;
  assign n17857 = ~n14045 & n17856;
  assign n17858 = ~n15657 & n17857;
  assign n17859 = ~n2543 & ~n3066;
  assign n17860 = ~n3983 & n17859;
  assign n17861 = ~n4024 & n17860;
  assign n17862 = ~n4999 & n17861;
  assign n17863 = ~n5827 & n17862;
  assign n17864 = ~n6893 & n17863;
  assign n17865 = ~n7890 & n17864;
  assign n17866 = ~n9131 & n17865;
  assign n17867 = ~n10278 & n17866;
  assign n17868 = ~n11662 & n17867;
  assign n17869 = ~n13191 & n17868;
  assign n17870 = ~n14848 & n17869;
  assign n17871 = ~n17858 & ~n17870;
  assign n17872 = n17854 & n17871;
  assign n17873 = n17838 & n17872;
  assign n17874 = n17806 & n17873;
  assign n17875 = n17773 & n17874;
  assign n17876 = ~n17749 & ~n17875;
  assign n17877 = ~n17738 & n17876;
  assign n17878 = pi028 & ~n16417;
  assign n17879 = ~n17766 & n17878;
  assign n17880 = ~n16216 & n17879;
  assign n17881 = ~n16215 & n17880;
  assign n17882 = n16222 & n17881;
  assign n17883 = n17637 & n17882;
  assign n17884 = n17629 & n17883;
  assign n17885 = n17765 & n17884;
  assign n17886 = n17874 & n17885;
  assign n17887 = ~n1739 & ~n9653;
  assign n17888 = n2317 & n17887;
  assign n17889 = n15961 & n17888;
  assign n17890 = ~pi263 & pi271;
  assign n17891 = pi265 & ~pi273;
  assign n17892 = ~pi265 & pi273;
  assign n17893 = pi266 & ~pi274;
  assign n17894 = ~pi266 & pi274;
  assign n17895 = pi267 & ~pi275;
  assign n17896 = ~pi267 & pi275;
  assign n17897 = pi268 & ~pi276;
  assign n17898 = ~pi268 & pi276;
  assign n17899 = ~pi269 & pi277;
  assign n17900 = pi270 & ~pi278;
  assign n17901 = ~n17899 & n17900;
  assign n17902 = pi269 & ~pi277;
  assign n17903 = ~n17901 & ~n17902;
  assign n17904 = ~n17898 & ~n17903;
  assign n17905 = ~n17897 & ~n17904;
  assign n17906 = ~n17896 & ~n17905;
  assign n17907 = ~n17895 & ~n17906;
  assign n17908 = ~n17894 & ~n17907;
  assign n17909 = ~n17893 & ~n17908;
  assign n17910 = ~n17892 & ~n17909;
  assign n17911 = ~n17891 & ~n17910;
  assign n17912 = pi264 & ~n17911;
  assign n17913 = ~pi264 & ~n17891;
  assign n17914 = ~n17910 & n17913;
  assign n17915 = ~pi272 & ~n17914;
  assign n17916 = pi263 & ~pi271;
  assign n17917 = ~n17915 & ~n17916;
  assign n17918 = ~n17912 & n17917;
  assign n17919 = ~n17890 & ~n17918;
  assign n17920 = n15960 & ~n17919;
  assign n17921 = n17889 & n17920;
  assign n17922 = n2316 & n14185;
  assign n17923 = ~n656 & ~n779;
  assign n17924 = n16011 & n17923;
  assign n17925 = n17922 & n17924;
  assign n17926 = ~n1432 & ~n1555;
  assign n17927 = n14181 & n17926;
  assign n17928 = n14421 & n17927;
  assign n17929 = n17925 & n17928;
  assign n17930 = ~n4429 & ~n4459;
  assign n17931 = n5732 & n17930;
  assign n17932 = ~n2542 & ~n3254;
  assign n17933 = n14137 & n17932;
  assign n17934 = n17931 & n17933;
  assign n17935 = ~n5626 & ~n5685;
  assign n17936 = n14144 & n17935;
  assign n17937 = n14142 & n17936;
  assign n17938 = n17934 & n17937;
  assign n17939 = ~n2423 & ~n2601;
  assign n17940 = n3819 & n17939;
  assign n17941 = ~n1404 & ~n1527;
  assign n17942 = n15966 & n17941;
  assign n17943 = n5716 & n17942;
  assign n17944 = ~n2484 & ~n2574;
  assign n17945 = n15964 & n17944;
  assign n17946 = n15970 & n17945;
  assign n17947 = n17943 & n17946;
  assign n17948 = ~n751 & ~n782;
  assign n17949 = n15978 & n17948;
  assign n17950 = pi029 & ~n501;
  assign n17951 = n12872 & n17950;
  assign n17952 = n17949 & n17951;
  assign n17953 = n12562 & n14191;
  assign n17954 = n5752 & n17953;
  assign n17955 = n17952 & n17954;
  assign n17956 = n17947 & n17955;
  assign n17957 = ~n14352 & ~n15989;
  assign n17958 = ~n16146 & n17957;
  assign n17959 = ~n8427 & ~n14387;
  assign n17960 = n15988 & n17959;
  assign n17961 = n15992 & n17960;
  assign n17962 = n17958 & n17961;
  assign n17963 = n7241 & n12544;
  assign n17964 = ~n5350 & ~n5658;
  assign n17965 = ~n5261 & ~n5599;
  assign n17966 = n17964 & n17965;
  assign n17967 = n17963 & n17966;
  assign n17968 = ~n7387 & ~n7477;
  assign n17969 = n16376 & n17968;
  assign n17970 = ~n6285 & ~n7664;
  assign n17971 = n16386 & n17970;
  assign n17972 = n17969 & n17971;
  assign n17973 = n17967 & n17972;
  assign n17974 = ~n3285 & ~n3622;
  assign n17975 = n4796 & n17974;
  assign n17976 = n14275 & n17975;
  assign n17977 = ~n4432 & ~n4580;
  assign n17978 = n5720 & n17977;
  assign n17979 = n15997 & n17978;
  assign n17980 = n17976 & n17979;
  assign n17981 = n17973 & n17980;
  assign n17982 = n17962 & n17981;
  assign n17983 = n17956 & n17982;
  assign n17984 = ~n1172 & n17983;
  assign n17985 = ~n996 & n17984;
  assign n17986 = ~n2306 & n17985;
  assign n17987 = ~n500 & n17986;
  assign n17988 = n17940 & n17987;
  assign n17989 = ~n3590 & ~n3649;
  assign n17990 = n14136 & n17989;
  assign n17991 = n14139 & n17990;
  assign n17992 = n17988 & n17991;
  assign n17993 = n17938 & n17992;
  assign n17994 = n17929 & n17993;
  assign n17995 = n17921 & n17994;
  assign n17996 = ~n14380 & ~n14415;
  assign n17997 = ~n15949 & ~n16174;
  assign n17998 = n17996 & n17997;
  assign n17999 = ~n12710 & ~n12772;
  assign n18000 = ~n12712 & ~n14176;
  assign n18001 = n17999 & n18000;
  assign n18002 = ~n11132 & ~n12808;
  assign n18003 = ~n12770 & ~n12810;
  assign n18004 = n18002 & n18003;
  assign n18005 = n18001 & n18004;
  assign n18006 = n17998 & n18005;
  assign n18007 = ~n9910 & n14131;
  assign n18008 = ~n9821 & ~n9912;
  assign n18009 = n18007 & n18008;
  assign n18010 = ~n6312 & ~n6341;
  assign n18011 = n6181 & n18010;
  assign n18012 = n16020 & n18011;
  assign n18013 = ~n7414 & ~n7750;
  assign n18014 = ~n8454 & ~n8483;
  assign n18015 = n18013 & n18014;
  assign n18016 = ~n7355 & ~n7504;
  assign n18017 = n8878 & n18016;
  assign n18018 = n18015 & n18017;
  assign n18019 = n18012 & n18018;
  assign n18020 = n18009 & n18019;
  assign n18021 = ~n11041 & ~n11069;
  assign n18022 = ~n11071 & ~n11130;
  assign n18023 = n18021 & n18022;
  assign n18024 = ~n9823 & ~n9851;
  assign n18025 = ~n9853 & ~n11039;
  assign n18026 = n18024 & n18025;
  assign n18027 = n18023 & n18026;
  assign n18028 = n18020 & n18027;
  assign n18029 = n18006 & n18028;
  assign n18030 = n17995 & n18029;
  assign n18031 = ~n6131 & n18030;
  assign n18032 = ~n1432 & ~n1525;
  assign n18033 = n14181 & n18032;
  assign n18034 = n17888 & n18033;
  assign n18035 = n15962 & n18034;
  assign n18036 = ~n1207 & ~n1237;
  assign n18037 = n12582 & n18036;
  assign n18038 = n3819 & n14143;
  assign n18039 = ~n1435 & ~n2147;
  assign n18040 = n15964 & n18039;
  assign n18041 = ~n1497 & ~n2082;
  assign n18042 = n15966 & n18041;
  assign n18043 = n18040 & n18042;
  assign n18044 = ~n2755 & ~n3682;
  assign n18045 = n14210 & n18044;
  assign n18046 = n12604 & n18045;
  assign n18047 = n18043 & n18046;
  assign n18048 = ~n659 & ~n1179;
  assign n18049 = n15978 & n18048;
  assign n18050 = pi030 & ~n501;
  assign n18051 = n12872 & n18050;
  assign n18052 = n18049 & n18051;
  assign n18053 = n12618 & n14253;
  assign n18054 = n18052 & n18053;
  assign n18055 = n18047 & n18054;
  assign n18056 = ~n14321 & ~n15989;
  assign n18057 = ~n16115 & ~n17890;
  assign n18058 = n18056 & n18057;
  assign n18059 = ~n8605 & ~n14387;
  assign n18060 = n15988 & n18059;
  assign n18061 = n15992 & n18060;
  assign n18062 = n18058 & n18061;
  assign n18063 = ~n6373 & ~n6615;
  assign n18064 = n7241 & n18063;
  assign n18065 = ~n5321 & ~n5350;
  assign n18066 = ~n4679 & ~n5599;
  assign n18067 = n18065 & n18066;
  assign n18068 = n18064 & n18067;
  assign n18069 = ~n7328 & ~n7635;
  assign n18070 = n16377 & n18069;
  assign n18071 = n14202 & n18070;
  assign n18072 = n18068 & n18071;
  assign n18073 = n12550 & n15998;
  assign n18074 = n15970 & n18073;
  assign n18075 = ~n4373 & ~n4402;
  assign n18076 = n5720 & n18075;
  assign n18077 = n11402 & n18076;
  assign n18078 = n18074 & n18077;
  assign n18079 = n18072 & n18078;
  assign n18080 = n18062 & n18079;
  assign n18081 = n18055 & n18080;
  assign n18082 = ~n1172 & n18081;
  assign n18083 = ~n996 & n18082;
  assign n18084 = ~n2306 & n18083;
  assign n18085 = ~n500 & n18084;
  assign n18086 = n18038 & n18085;
  assign n18087 = n18037 & n18086;
  assign n18088 = n14421 & n17922;
  assign n18089 = n18087 & n18088;
  assign n18090 = ~n5348 & ~n5377;
  assign n18091 = n16032 & n18090;
  assign n18092 = ~n4400 & ~n5597;
  assign n18093 = n16034 & n18092;
  assign n18094 = n18091 & n18093;
  assign n18095 = n16021 & n18094;
  assign n18096 = ~n3709 & ~n3738;
  assign n18097 = n16028 & n18096;
  assign n18098 = ~n2662 & ~n2782;
  assign n18099 = ~n2691 & ~n2721;
  assign n18100 = n18098 & n18099;
  assign n18101 = n18097 & n18100;
  assign n18102 = n5732 & n14141;
  assign n18103 = n14137 & n16026;
  assign n18104 = n18102 & n18103;
  assign n18105 = n18101 & n18104;
  assign n18106 = n18095 & n18105;
  assign n18107 = n18089 & n18106;
  assign n18108 = n18035 & n18107;
  assign n18109 = ~n15949 & ~n16143;
  assign n18110 = ~n17918 & n18109;
  assign n18111 = ~n14349 & ~n14415;
  assign n18112 = n18000 & n18111;
  assign n18113 = ~n12740 & ~n12810;
  assign n18114 = ~n12710 & ~n12742;
  assign n18115 = n18113 & n18114;
  assign n18116 = n18112 & n18115;
  assign n18117 = n18110 & n18116;
  assign n18118 = ~n9762 & ~n9821;
  assign n18119 = n18024 & n18118;
  assign n18120 = ~n8483 & ~n8632;
  assign n18121 = n10824 & n18120;
  assign n18122 = ~n6400 & ~n7662;
  assign n18123 = n14132 & n18122;
  assign n18124 = n18121 & n18123;
  assign n18125 = ~n9760 & n14131;
  assign n18126 = n18124 & n18125;
  assign n18127 = n18119 & n18126;
  assign n18128 = n18002 & n18022;
  assign n18129 = ~n9853 & ~n11165;
  assign n18130 = ~n11069 & ~n11167;
  assign n18131 = n18129 & n18130;
  assign n18132 = n18128 & n18131;
  assign n18133 = n18127 & n18132;
  assign n18134 = n18117 & n18133;
  assign n18135 = n18108 & n18134;
  assign n18136 = ~n6131 & n18135;
  assign n18137 = ~n18031 & ~n18136;
  assign n18138 = n16192 & ~n18137;
  assign n18139 = ~n8867 & n18138;
  assign n18140 = ~n7235 & n18139;
  assign n18141 = n7296 & n18140;
  assign n18142 = n7231 & n18141;
  assign n18143 = ~n10027 & n18142;
  assign n18144 = ~n8866 & n18143;
  assign n18145 = n8898 & n18144;
  assign n18146 = n8863 & n18145;
  assign n18147 = ~n10788 & n18146;
  assign n18148 = ~n10026 & n18147;
  assign n18149 = n10072 & n18148;
  assign n18150 = n10021 & n18149;
  assign n18151 = ~n17886 & ~n18150;
  assign po015 = n17877 | ~n18151;
  assign n18153 = pi047 & ~n501;
  assign n18154 = ~n500 & n18153;
  assign n18155 = pi039 & ~n1173;
  assign n18156 = ~n1144 & n18155;
  assign n18157 = ~n1115 & n18156;
  assign n18158 = ~n1086 & n18157;
  assign n18159 = n1057 & n18158;
  assign n18160 = n1239 & n18159;
  assign n18161 = n1360 & n18160;
  assign n18162 = n968 & n18161;
  assign n18163 = n845 & n18162;
  assign po024 = n18154 | n18163;
  assign n18165 = pi048 & ~n501;
  assign n18166 = ~n500 & n18165;
  assign n18167 = pi040 & ~n1173;
  assign n18168 = ~n1144 & n18167;
  assign n18169 = ~n1115 & n18168;
  assign n18170 = ~n1086 & n18169;
  assign n18171 = n1057 & n18170;
  assign n18172 = n1239 & n18171;
  assign n18173 = n1360 & n18172;
  assign n18174 = n968 & n18173;
  assign n18175 = n845 & n18174;
  assign po025 = n18166 | n18175;
  assign n18177 = pi049 & ~n501;
  assign n18178 = ~n500 & n18177;
  assign n18179 = pi041 & ~n1173;
  assign n18180 = ~n1144 & n18179;
  assign n18181 = ~n1115 & n18180;
  assign n18182 = ~n1086 & n18181;
  assign n18183 = n1057 & n18182;
  assign n18184 = n1239 & n18183;
  assign n18185 = n1360 & n18184;
  assign n18186 = n968 & n18185;
  assign n18187 = n845 & n18186;
  assign po026 = n18178 | n18187;
  assign n18189 = pi050 & ~n501;
  assign n18190 = ~n500 & n18189;
  assign n18191 = pi042 & ~n1173;
  assign n18192 = ~n1144 & n18191;
  assign n18193 = ~n1115 & n18192;
  assign n18194 = ~n1086 & n18193;
  assign n18195 = n1057 & n18194;
  assign n18196 = n1239 & n18195;
  assign n18197 = n1360 & n18196;
  assign n18198 = n968 & n18197;
  assign n18199 = n845 & n18198;
  assign po027 = n18190 | n18199;
  assign n18201 = pi051 & ~n501;
  assign n18202 = ~n500 & n18201;
  assign n18203 = pi043 & ~n1173;
  assign n18204 = ~n1144 & n18203;
  assign n18205 = ~n1115 & n18204;
  assign n18206 = ~n1086 & n18205;
  assign n18207 = n1057 & n18206;
  assign n18208 = n1239 & n18207;
  assign n18209 = n1360 & n18208;
  assign n18210 = n968 & n18209;
  assign n18211 = n845 & n18210;
  assign po028 = n18202 | n18211;
  assign n18213 = pi052 & ~n501;
  assign n18214 = ~n500 & n18213;
  assign n18215 = pi044 & ~n1173;
  assign n18216 = ~n1144 & n18215;
  assign n18217 = ~n1115 & n18216;
  assign n18218 = ~n1086 & n18217;
  assign n18219 = n1057 & n18218;
  assign n18220 = n1239 & n18219;
  assign n18221 = n1360 & n18220;
  assign n18222 = n968 & n18221;
  assign n18223 = n845 & n18222;
  assign po029 = n18214 | n18223;
  assign n18225 = pi053 & ~n501;
  assign n18226 = ~n500 & n18225;
  assign n18227 = pi045 & ~n1173;
  assign n18228 = ~n1144 & n18227;
  assign n18229 = ~n1115 & n18228;
  assign n18230 = ~n1086 & n18229;
  assign n18231 = n1057 & n18230;
  assign n18232 = n1239 & n18231;
  assign n18233 = n1360 & n18232;
  assign n18234 = n968 & n18233;
  assign n18235 = n845 & n18234;
  assign po030 = n18226 | n18235;
  assign n18237 = pi054 & ~n501;
  assign n18238 = ~n500 & n18237;
  assign n18239 = pi046 & ~n1173;
  assign n18240 = ~n1144 & n18239;
  assign n18241 = ~n1115 & n18240;
  assign n18242 = ~n1086 & n18241;
  assign n18243 = n1057 & n18242;
  assign n18244 = n1239 & n18243;
  assign n18245 = n1360 & n18244;
  assign n18246 = n968 & n18245;
  assign n18247 = n845 & n18246;
  assign po031 = n18238 | n18247;
  assign n18249 = pi055 & ~n501;
  assign n18250 = ~n500 & n18249;
  assign n18251 = ~n2143 & n18250;
  assign n18252 = n2207 & n18251;
  assign n18253 = n2113 & n18252;
  assign n18254 = n1990 & n18253;
  assign n18255 = n1867 & n18254;
  assign n18256 = n1744 & n18255;
  assign n18257 = ~n1373 & n18256;
  assign n18258 = n2215 & n18162;
  assign n18259 = ~n1372 & n18258;
  assign n18260 = pi063 & ~n501;
  assign n18261 = n2219 & n18260;
  assign n18262 = ~n500 & n18261;
  assign n18263 = n2222 & n18262;
  assign n18264 = pi047 & ~n1173;
  assign n18265 = ~n1144 & n18264;
  assign n18266 = ~n1115 & n18265;
  assign n18267 = ~n1086 & n18266;
  assign n18268 = n1057 & n18267;
  assign n18269 = n1239 & n18268;
  assign n18270 = n1360 & n18269;
  assign n18271 = n968 & n18270;
  assign n18272 = n845 & n18271;
  assign n18273 = ~n18263 & ~n18272;
  assign n18274 = ~n18259 & n18273;
  assign po032 = n18257 | ~n18274;
  assign n18276 = pi056 & ~n501;
  assign n18277 = ~n500 & n18276;
  assign n18278 = ~n2143 & n18277;
  assign n18279 = n2207 & n18278;
  assign n18280 = n2113 & n18279;
  assign n18281 = n1990 & n18280;
  assign n18282 = n1867 & n18281;
  assign n18283 = n1744 & n18282;
  assign n18284 = ~n1373 & n18283;
  assign n18285 = n2215 & n18174;
  assign n18286 = ~n1372 & n18285;
  assign n18287 = pi064 & ~n501;
  assign n18288 = n2219 & n18287;
  assign n18289 = ~n500 & n18288;
  assign n18290 = n2222 & n18289;
  assign n18291 = pi048 & ~n1173;
  assign n18292 = ~n1144 & n18291;
  assign n18293 = ~n1115 & n18292;
  assign n18294 = ~n1086 & n18293;
  assign n18295 = n1057 & n18294;
  assign n18296 = n1239 & n18295;
  assign n18297 = n1360 & n18296;
  assign n18298 = n968 & n18297;
  assign n18299 = n845 & n18298;
  assign n18300 = ~n18290 & ~n18299;
  assign n18301 = ~n18286 & n18300;
  assign po033 = n18284 | ~n18301;
  assign n18303 = pi057 & ~n501;
  assign n18304 = ~n500 & n18303;
  assign n18305 = ~n2143 & n18304;
  assign n18306 = n2207 & n18305;
  assign n18307 = n2113 & n18306;
  assign n18308 = n1990 & n18307;
  assign n18309 = n1867 & n18308;
  assign n18310 = n1744 & n18309;
  assign n18311 = ~n1373 & n18310;
  assign n18312 = n2215 & n18186;
  assign n18313 = ~n1372 & n18312;
  assign n18314 = pi065 & ~n501;
  assign n18315 = n2219 & n18314;
  assign n18316 = ~n500 & n18315;
  assign n18317 = n2222 & n18316;
  assign n18318 = pi049 & ~n1173;
  assign n18319 = ~n1144 & n18318;
  assign n18320 = ~n1115 & n18319;
  assign n18321 = ~n1086 & n18320;
  assign n18322 = n1057 & n18321;
  assign n18323 = n1239 & n18322;
  assign n18324 = n1360 & n18323;
  assign n18325 = n968 & n18324;
  assign n18326 = n845 & n18325;
  assign n18327 = ~n18317 & ~n18326;
  assign n18328 = ~n18313 & n18327;
  assign po034 = n18311 | ~n18328;
  assign n18330 = pi058 & ~n501;
  assign n18331 = ~n500 & n18330;
  assign n18332 = ~n2143 & n18331;
  assign n18333 = n2207 & n18332;
  assign n18334 = n2113 & n18333;
  assign n18335 = n1990 & n18334;
  assign n18336 = n1867 & n18335;
  assign n18337 = n1744 & n18336;
  assign n18338 = ~n1373 & n18337;
  assign n18339 = n2215 & n18198;
  assign n18340 = ~n1372 & n18339;
  assign n18341 = pi066 & ~n501;
  assign n18342 = n2219 & n18341;
  assign n18343 = ~n500 & n18342;
  assign n18344 = n2222 & n18343;
  assign n18345 = pi050 & ~n1173;
  assign n18346 = ~n1144 & n18345;
  assign n18347 = ~n1115 & n18346;
  assign n18348 = ~n1086 & n18347;
  assign n18349 = n1057 & n18348;
  assign n18350 = n1239 & n18349;
  assign n18351 = n1360 & n18350;
  assign n18352 = n968 & n18351;
  assign n18353 = n845 & n18352;
  assign n18354 = ~n18344 & ~n18353;
  assign n18355 = ~n18340 & n18354;
  assign po035 = n18338 | ~n18355;
  assign n18357 = pi059 & ~n501;
  assign n18358 = ~n500 & n18357;
  assign n18359 = ~n2143 & n18358;
  assign n18360 = n2207 & n18359;
  assign n18361 = n2113 & n18360;
  assign n18362 = n1990 & n18361;
  assign n18363 = n1867 & n18362;
  assign n18364 = n1744 & n18363;
  assign n18365 = ~n1373 & n18364;
  assign n18366 = n2215 & n18210;
  assign n18367 = ~n1372 & n18366;
  assign n18368 = pi067 & ~n501;
  assign n18369 = n2219 & n18368;
  assign n18370 = ~n500 & n18369;
  assign n18371 = n2222 & n18370;
  assign n18372 = pi051 & ~n1173;
  assign n18373 = ~n1144 & n18372;
  assign n18374 = ~n1115 & n18373;
  assign n18375 = ~n1086 & n18374;
  assign n18376 = n1057 & n18375;
  assign n18377 = n1239 & n18376;
  assign n18378 = n1360 & n18377;
  assign n18379 = n968 & n18378;
  assign n18380 = n845 & n18379;
  assign n18381 = ~n18371 & ~n18380;
  assign n18382 = ~n18367 & n18381;
  assign po036 = n18365 | ~n18382;
  assign n18384 = pi060 & ~n501;
  assign n18385 = ~n500 & n18384;
  assign n18386 = ~n2143 & n18385;
  assign n18387 = n2207 & n18386;
  assign n18388 = n2113 & n18387;
  assign n18389 = n1990 & n18388;
  assign n18390 = n1867 & n18389;
  assign n18391 = n1744 & n18390;
  assign n18392 = ~n1373 & n18391;
  assign n18393 = n2215 & n18222;
  assign n18394 = ~n1372 & n18393;
  assign n18395 = pi068 & ~n501;
  assign n18396 = n2219 & n18395;
  assign n18397 = ~n500 & n18396;
  assign n18398 = n2222 & n18397;
  assign n18399 = pi052 & ~n1173;
  assign n18400 = ~n1144 & n18399;
  assign n18401 = ~n1115 & n18400;
  assign n18402 = ~n1086 & n18401;
  assign n18403 = n1057 & n18402;
  assign n18404 = n1239 & n18403;
  assign n18405 = n1360 & n18404;
  assign n18406 = n968 & n18405;
  assign n18407 = n845 & n18406;
  assign n18408 = ~n18398 & ~n18407;
  assign n18409 = ~n18394 & n18408;
  assign po037 = n18392 | ~n18409;
  assign n18411 = pi061 & ~n501;
  assign n18412 = ~n500 & n18411;
  assign n18413 = ~n2143 & n18412;
  assign n18414 = n2207 & n18413;
  assign n18415 = n2113 & n18414;
  assign n18416 = n1990 & n18415;
  assign n18417 = n1867 & n18416;
  assign n18418 = n1744 & n18417;
  assign n18419 = ~n1373 & n18418;
  assign n18420 = n2215 & n18234;
  assign n18421 = ~n1372 & n18420;
  assign n18422 = pi069 & ~n501;
  assign n18423 = n2219 & n18422;
  assign n18424 = ~n500 & n18423;
  assign n18425 = n2222 & n18424;
  assign n18426 = pi053 & ~n1173;
  assign n18427 = ~n1144 & n18426;
  assign n18428 = ~n1115 & n18427;
  assign n18429 = ~n1086 & n18428;
  assign n18430 = n1057 & n18429;
  assign n18431 = n1239 & n18430;
  assign n18432 = n1360 & n18431;
  assign n18433 = n968 & n18432;
  assign n18434 = n845 & n18433;
  assign n18435 = ~n18425 & ~n18434;
  assign n18436 = ~n18421 & n18435;
  assign po038 = n18419 | ~n18436;
  assign n18438 = pi062 & ~n501;
  assign n18439 = ~n500 & n18438;
  assign n18440 = ~n2143 & n18439;
  assign n18441 = n2207 & n18440;
  assign n18442 = n2113 & n18441;
  assign n18443 = n1990 & n18442;
  assign n18444 = n1867 & n18443;
  assign n18445 = n1744 & n18444;
  assign n18446 = ~n1373 & n18445;
  assign n18447 = n2215 & n18246;
  assign n18448 = ~n1372 & n18447;
  assign n18449 = pi070 & ~n501;
  assign n18450 = n2219 & n18449;
  assign n18451 = ~n500 & n18450;
  assign n18452 = n2222 & n18451;
  assign n18453 = pi054 & ~n1173;
  assign n18454 = ~n1144 & n18453;
  assign n18455 = ~n1115 & n18454;
  assign n18456 = ~n1086 & n18455;
  assign n18457 = n1057 & n18456;
  assign n18458 = n1239 & n18457;
  assign n18459 = n1360 & n18458;
  assign n18460 = n968 & n18459;
  assign n18461 = n845 & n18460;
  assign n18462 = ~n18452 & ~n18461;
  assign n18463 = ~n18448 & n18462;
  assign po039 = n18446 | ~n18463;
  assign n18465 = pi055 & ~n2143;
  assign n18466 = n2207 & n18465;
  assign n18467 = n2113 & n18466;
  assign n18468 = n1990 & n18467;
  assign n18469 = n1867 & n18468;
  assign n18470 = n2253 & n18469;
  assign n18471 = ~n2245 & n18470;
  assign n18472 = ~n2244 & n18471;
  assign n18473 = ~n2242 & n18472;
  assign n18474 = n1359 & n18159;
  assign n18475 = n2272 & n18474;
  assign n18476 = n2271 & n18475;
  assign n18477 = n2268 & n18476;
  assign n18478 = ~n1372 & n18477;
  assign n18479 = ~n2243 & n18478;
  assign n18480 = ~n2263 & n18479;
  assign n18481 = pi079 & ~n501;
  assign n18482 = n2311 & n18481;
  assign n18483 = n2309 & n18482;
  assign n18484 = ~n2306 & n18483;
  assign n18485 = ~n500 & n18484;
  assign n18486 = n2318 & n18485;
  assign n18487 = ~n18480 & ~n18486;
  assign n18488 = ~n18473 & n18487;
  assign n18489 = pi063 & ~po145;
  assign n18490 = ~n2245 & n18489;
  assign n18491 = ~n2324 & n18490;
  assign n18492 = ~n2322 & n18491;
  assign n18493 = pi071 & ~n501;
  assign n18494 = n2219 & n18493;
  assign n18495 = ~n500 & n18494;
  assign n18496 = n2394 & n18495;
  assign n18497 = n2846 & n18496;
  assign n18498 = n3056 & n18497;
  assign n18499 = ~n2331 & n18498;
  assign n18500 = ~n2329 & n18499;
  assign n18501 = ~n18492 & ~n18500;
  assign po040 = ~n18488 | ~n18501;
  assign n18503 = pi056 & ~n2143;
  assign n18504 = n2207 & n18503;
  assign n18505 = n2113 & n18504;
  assign n18506 = n1990 & n18505;
  assign n18507 = n1867 & n18506;
  assign n18508 = n2253 & n18507;
  assign n18509 = ~n2245 & n18508;
  assign n18510 = ~n2244 & n18509;
  assign n18511 = ~n2242 & n18510;
  assign n18512 = n1359 & n18171;
  assign n18513 = n2272 & n18512;
  assign n18514 = n2271 & n18513;
  assign n18515 = n2268 & n18514;
  assign n18516 = ~n1372 & n18515;
  assign n18517 = ~n2243 & n18516;
  assign n18518 = ~n2263 & n18517;
  assign n18519 = pi080 & ~n501;
  assign n18520 = n2311 & n18519;
  assign n18521 = n2309 & n18520;
  assign n18522 = ~n2306 & n18521;
  assign n18523 = ~n500 & n18522;
  assign n18524 = n2318 & n18523;
  assign n18525 = ~n18518 & ~n18524;
  assign n18526 = ~n18511 & n18525;
  assign n18527 = pi064 & ~po145;
  assign n18528 = ~n2245 & n18527;
  assign n18529 = ~n2324 & n18528;
  assign n18530 = ~n2322 & n18529;
  assign n18531 = pi072 & ~n501;
  assign n18532 = n2219 & n18531;
  assign n18533 = ~n500 & n18532;
  assign n18534 = n2394 & n18533;
  assign n18535 = n2846 & n18534;
  assign n18536 = n3056 & n18535;
  assign n18537 = ~n2331 & n18536;
  assign n18538 = ~n2329 & n18537;
  assign n18539 = ~n18530 & ~n18538;
  assign po041 = ~n18526 | ~n18539;
  assign n18541 = pi057 & ~n2143;
  assign n18542 = n2207 & n18541;
  assign n18543 = n2113 & n18542;
  assign n18544 = n1990 & n18543;
  assign n18545 = n1867 & n18544;
  assign n18546 = n2253 & n18545;
  assign n18547 = ~n2245 & n18546;
  assign n18548 = ~n2244 & n18547;
  assign n18549 = ~n2242 & n18548;
  assign n18550 = n1359 & n18183;
  assign n18551 = n2272 & n18550;
  assign n18552 = n2271 & n18551;
  assign n18553 = n2268 & n18552;
  assign n18554 = ~n1372 & n18553;
  assign n18555 = ~n2243 & n18554;
  assign n18556 = ~n2263 & n18555;
  assign n18557 = pi081 & ~n501;
  assign n18558 = n2311 & n18557;
  assign n18559 = n2309 & n18558;
  assign n18560 = ~n2306 & n18559;
  assign n18561 = ~n500 & n18560;
  assign n18562 = n2318 & n18561;
  assign n18563 = ~n18556 & ~n18562;
  assign n18564 = ~n18549 & n18563;
  assign n18565 = pi065 & ~po145;
  assign n18566 = ~n2245 & n18565;
  assign n18567 = ~n2324 & n18566;
  assign n18568 = ~n2322 & n18567;
  assign n18569 = pi073 & ~n501;
  assign n18570 = n2219 & n18569;
  assign n18571 = ~n500 & n18570;
  assign n18572 = n2394 & n18571;
  assign n18573 = n2846 & n18572;
  assign n18574 = n3056 & n18573;
  assign n18575 = ~n2331 & n18574;
  assign n18576 = ~n2329 & n18575;
  assign n18577 = ~n18568 & ~n18576;
  assign po042 = ~n18564 | ~n18577;
  assign n18579 = pi058 & ~n2143;
  assign n18580 = n2207 & n18579;
  assign n18581 = n2113 & n18580;
  assign n18582 = n1990 & n18581;
  assign n18583 = n1867 & n18582;
  assign n18584 = n2253 & n18583;
  assign n18585 = ~n2245 & n18584;
  assign n18586 = ~n2244 & n18585;
  assign n18587 = ~n2242 & n18586;
  assign n18588 = n1359 & n18195;
  assign n18589 = n2272 & n18588;
  assign n18590 = n2271 & n18589;
  assign n18591 = n2268 & n18590;
  assign n18592 = ~n1372 & n18591;
  assign n18593 = ~n2243 & n18592;
  assign n18594 = ~n2263 & n18593;
  assign n18595 = pi082 & ~n501;
  assign n18596 = n2311 & n18595;
  assign n18597 = n2309 & n18596;
  assign n18598 = ~n2306 & n18597;
  assign n18599 = ~n500 & n18598;
  assign n18600 = n2318 & n18599;
  assign n18601 = ~n18594 & ~n18600;
  assign n18602 = ~n18587 & n18601;
  assign n18603 = pi066 & ~po145;
  assign n18604 = ~n2245 & n18603;
  assign n18605 = ~n2324 & n18604;
  assign n18606 = ~n2322 & n18605;
  assign n18607 = pi074 & ~n501;
  assign n18608 = n2219 & n18607;
  assign n18609 = ~n500 & n18608;
  assign n18610 = n2394 & n18609;
  assign n18611 = n2846 & n18610;
  assign n18612 = n3056 & n18611;
  assign n18613 = ~n2331 & n18612;
  assign n18614 = ~n2329 & n18613;
  assign n18615 = ~n18606 & ~n18614;
  assign po043 = ~n18602 | ~n18615;
  assign n18617 = pi059 & ~n2143;
  assign n18618 = n2207 & n18617;
  assign n18619 = n2113 & n18618;
  assign n18620 = n1990 & n18619;
  assign n18621 = n1867 & n18620;
  assign n18622 = n2253 & n18621;
  assign n18623 = ~n2245 & n18622;
  assign n18624 = ~n2244 & n18623;
  assign n18625 = ~n2242 & n18624;
  assign n18626 = n1359 & n18207;
  assign n18627 = n2272 & n18626;
  assign n18628 = n2271 & n18627;
  assign n18629 = n2268 & n18628;
  assign n18630 = ~n1372 & n18629;
  assign n18631 = ~n2243 & n18630;
  assign n18632 = ~n2263 & n18631;
  assign n18633 = pi083 & ~n501;
  assign n18634 = n2311 & n18633;
  assign n18635 = n2309 & n18634;
  assign n18636 = ~n2306 & n18635;
  assign n18637 = ~n500 & n18636;
  assign n18638 = n2318 & n18637;
  assign n18639 = ~n18632 & ~n18638;
  assign n18640 = ~n18625 & n18639;
  assign n18641 = pi067 & ~po145;
  assign n18642 = ~n2245 & n18641;
  assign n18643 = ~n2324 & n18642;
  assign n18644 = ~n2322 & n18643;
  assign n18645 = pi075 & ~n501;
  assign n18646 = n2219 & n18645;
  assign n18647 = ~n500 & n18646;
  assign n18648 = n2394 & n18647;
  assign n18649 = n2846 & n18648;
  assign n18650 = n3056 & n18649;
  assign n18651 = ~n2331 & n18650;
  assign n18652 = ~n2329 & n18651;
  assign n18653 = ~n18644 & ~n18652;
  assign po044 = ~n18640 | ~n18653;
  assign n18655 = pi060 & ~n2143;
  assign n18656 = n2207 & n18655;
  assign n18657 = n2113 & n18656;
  assign n18658 = n1990 & n18657;
  assign n18659 = n1867 & n18658;
  assign n18660 = n2253 & n18659;
  assign n18661 = ~n2245 & n18660;
  assign n18662 = ~n2244 & n18661;
  assign n18663 = ~n2242 & n18662;
  assign n18664 = n1359 & n18219;
  assign n18665 = n2272 & n18664;
  assign n18666 = n2271 & n18665;
  assign n18667 = n2268 & n18666;
  assign n18668 = ~n1372 & n18667;
  assign n18669 = ~n2243 & n18668;
  assign n18670 = ~n2263 & n18669;
  assign n18671 = pi084 & ~n501;
  assign n18672 = n2311 & n18671;
  assign n18673 = n2309 & n18672;
  assign n18674 = ~n2306 & n18673;
  assign n18675 = ~n500 & n18674;
  assign n18676 = n2318 & n18675;
  assign n18677 = ~n18670 & ~n18676;
  assign n18678 = ~n18663 & n18677;
  assign n18679 = pi068 & ~po145;
  assign n18680 = ~n2245 & n18679;
  assign n18681 = ~n2324 & n18680;
  assign n18682 = ~n2322 & n18681;
  assign n18683 = pi076 & ~n501;
  assign n18684 = n2219 & n18683;
  assign n18685 = ~n500 & n18684;
  assign n18686 = n2394 & n18685;
  assign n18687 = n2846 & n18686;
  assign n18688 = n3056 & n18687;
  assign n18689 = ~n2331 & n18688;
  assign n18690 = ~n2329 & n18689;
  assign n18691 = ~n18682 & ~n18690;
  assign po045 = ~n18678 | ~n18691;
  assign n18693 = pi061 & ~n2143;
  assign n18694 = n2207 & n18693;
  assign n18695 = n2113 & n18694;
  assign n18696 = n1990 & n18695;
  assign n18697 = n1867 & n18696;
  assign n18698 = n2253 & n18697;
  assign n18699 = ~n2245 & n18698;
  assign n18700 = ~n2244 & n18699;
  assign n18701 = ~n2242 & n18700;
  assign n18702 = n1359 & n18231;
  assign n18703 = n2272 & n18702;
  assign n18704 = n2271 & n18703;
  assign n18705 = n2268 & n18704;
  assign n18706 = ~n1372 & n18705;
  assign n18707 = ~n2243 & n18706;
  assign n18708 = ~n2263 & n18707;
  assign n18709 = pi085 & ~n501;
  assign n18710 = n2311 & n18709;
  assign n18711 = n2309 & n18710;
  assign n18712 = ~n2306 & n18711;
  assign n18713 = ~n500 & n18712;
  assign n18714 = n2318 & n18713;
  assign n18715 = ~n18708 & ~n18714;
  assign n18716 = ~n18701 & n18715;
  assign n18717 = pi069 & ~po145;
  assign n18718 = ~n2245 & n18717;
  assign n18719 = ~n2324 & n18718;
  assign n18720 = ~n2322 & n18719;
  assign n18721 = pi077 & ~n501;
  assign n18722 = n2219 & n18721;
  assign n18723 = ~n500 & n18722;
  assign n18724 = n2394 & n18723;
  assign n18725 = n2846 & n18724;
  assign n18726 = n3056 & n18725;
  assign n18727 = ~n2331 & n18726;
  assign n18728 = ~n2329 & n18727;
  assign n18729 = ~n18720 & ~n18728;
  assign po046 = ~n18716 | ~n18729;
  assign n18731 = pi062 & ~n2143;
  assign n18732 = n2207 & n18731;
  assign n18733 = n2113 & n18732;
  assign n18734 = n1990 & n18733;
  assign n18735 = n1867 & n18734;
  assign n18736 = n2253 & n18735;
  assign n18737 = ~n2245 & n18736;
  assign n18738 = ~n2244 & n18737;
  assign n18739 = ~n2242 & n18738;
  assign n18740 = n1359 & n18243;
  assign n18741 = n2272 & n18740;
  assign n18742 = n2271 & n18741;
  assign n18743 = n2268 & n18742;
  assign n18744 = ~n1372 & n18743;
  assign n18745 = ~n2243 & n18744;
  assign n18746 = ~n2263 & n18745;
  assign n18747 = pi086 & ~n501;
  assign n18748 = n2311 & n18747;
  assign n18749 = n2309 & n18748;
  assign n18750 = ~n2306 & n18749;
  assign n18751 = ~n500 & n18750;
  assign n18752 = n2318 & n18751;
  assign n18753 = ~n18746 & ~n18752;
  assign n18754 = ~n18739 & n18753;
  assign n18755 = pi070 & ~po145;
  assign n18756 = ~n2245 & n18755;
  assign n18757 = ~n2324 & n18756;
  assign n18758 = ~n2322 & n18757;
  assign n18759 = pi078 & ~n501;
  assign n18760 = n2219 & n18759;
  assign n18761 = ~n500 & n18760;
  assign n18762 = n2394 & n18761;
  assign n18763 = n2846 & n18762;
  assign n18764 = n3056 & n18763;
  assign n18765 = ~n2331 & n18764;
  assign n18766 = ~n2329 & n18765;
  assign n18767 = ~n18758 & ~n18766;
  assign po047 = ~n18754 | ~n18767;
  assign n18769 = pi087 & ~n501;
  assign n18770 = n2311 & n18769;
  assign n18771 = n2309 & n18770;
  assign n18772 = ~n2306 & n18771;
  assign n18773 = ~n500 & n18772;
  assign n18774 = n2316 & n18773;
  assign n18775 = n3555 & n18774;
  assign n18776 = n3801 & n18775;
  assign n18777 = n3495 & n18776;
  assign n18778 = n3226 & n18777;
  assign n18779 = ~n3107 & n18778;
  assign n18780 = ~n3097 & n18779;
  assign n18781 = ~n3067 & n18780;
  assign n18782 = ~n3828 & n18489;
  assign n18783 = n3833 & n18782;
  assign n18784 = pi095 & ~n501;
  assign n18785 = n2311 & n18784;
  assign n18786 = n3813 & n18785;
  assign n18787 = n3811 & n18786;
  assign n18788 = ~n2306 & n18787;
  assign n18789 = n3819 & n18788;
  assign n18790 = n3823 & n18789;
  assign n18791 = n3809 & n18790;
  assign n18792 = ~n18783 & ~n18791;
  assign n18793 = ~n18781 & n18792;
  assign n18794 = pi071 & ~n2363;
  assign n18795 = n3847 & n18794;
  assign n18796 = n3855 & n18795;
  assign n18797 = n3843 & n18796;
  assign n18798 = n3869 & n18797;
  assign n18799 = ~n3066 & n18798;
  assign n18800 = n3874 & n18799;
  assign n18801 = ~n3837 & n18800;
  assign n18802 = ~n1897 & n18465;
  assign n18803 = n3082 & n18802;
  assign n18804 = n3888 & n18803;
  assign n18805 = ~n3886 & n18804;
  assign n18806 = n3885 & n18805;
  assign n18807 = ~n2242 & n18806;
  assign n18808 = ~n3095 & n18807;
  assign n18809 = ~n3878 & n18808;
  assign n18810 = ~n3877 & n18809;
  assign n18811 = ~n3837 & n18810;
  assign n18812 = ~n18801 & ~n18811;
  assign n18813 = pi079 & ~n3864;
  assign n18814 = ~n3919 & n18813;
  assign n18815 = ~n3916 & n18814;
  assign n18816 = n3924 & n18815;
  assign n18817 = n3903 & n18475;
  assign n18818 = n3907 & n18817;
  assign n18819 = ~n1372 & n18818;
  assign n18820 = ~n2243 & n18819;
  assign n18821 = ~n3104 & n18820;
  assign n18822 = ~n3901 & n18821;
  assign n18823 = ~n3837 & n18822;
  assign n18824 = ~n3900 & n18823;
  assign n18825 = ~n18816 & ~n18824;
  assign n18826 = n18812 & n18825;
  assign po048 = ~n18793 | ~n18826;
  assign n18828 = pi072 & ~n2363;
  assign n18829 = n3847 & n18828;
  assign n18830 = n3855 & n18829;
  assign n18831 = n3843 & n18830;
  assign n18832 = n3869 & n18831;
  assign n18833 = ~n3066 & n18832;
  assign n18834 = n3874 & n18833;
  assign n18835 = ~n3837 & n18834;
  assign n18836 = ~n3828 & n18527;
  assign n18837 = n3833 & n18836;
  assign n18838 = pi096 & ~n501;
  assign n18839 = n2311 & n18838;
  assign n18840 = n3813 & n18839;
  assign n18841 = n3811 & n18840;
  assign n18842 = ~n2306 & n18841;
  assign n18843 = n3819 & n18842;
  assign n18844 = n3823 & n18843;
  assign n18845 = n3809 & n18844;
  assign n18846 = ~n18837 & ~n18845;
  assign n18847 = ~n18835 & n18846;
  assign n18848 = pi088 & ~n501;
  assign n18849 = n2311 & n18848;
  assign n18850 = n2309 & n18849;
  assign n18851 = ~n2306 & n18850;
  assign n18852 = ~n500 & n18851;
  assign n18853 = n2316 & n18852;
  assign n18854 = n3555 & n18853;
  assign n18855 = n3801 & n18854;
  assign n18856 = n3495 & n18855;
  assign n18857 = n3226 & n18856;
  assign n18858 = ~n3107 & n18857;
  assign n18859 = ~n3097 & n18858;
  assign n18860 = ~n3067 & n18859;
  assign n18861 = ~n1897 & n18503;
  assign n18862 = n3082 & n18861;
  assign n18863 = n3888 & n18862;
  assign n18864 = ~n3886 & n18863;
  assign n18865 = n3885 & n18864;
  assign n18866 = ~n2242 & n18865;
  assign n18867 = ~n3095 & n18866;
  assign n18868 = ~n3878 & n18867;
  assign n18869 = ~n3877 & n18868;
  assign n18870 = ~n3837 & n18869;
  assign n18871 = ~n18860 & ~n18870;
  assign n18872 = n3903 & n18513;
  assign n18873 = n3907 & n18872;
  assign n18874 = ~n1372 & n18873;
  assign n18875 = ~n2243 & n18874;
  assign n18876 = ~n3104 & n18875;
  assign n18877 = ~n3901 & n18876;
  assign n18878 = ~n3837 & n18877;
  assign n18879 = ~n3900 & n18878;
  assign n18880 = pi080 & ~n3864;
  assign n18881 = ~n3919 & n18880;
  assign n18882 = ~n3916 & n18881;
  assign n18883 = n3924 & n18882;
  assign n18884 = ~n18879 & ~n18883;
  assign n18885 = n18871 & n18884;
  assign po049 = ~n18847 | ~n18885;
  assign n18887 = pi089 & ~n501;
  assign n18888 = n2311 & n18887;
  assign n18889 = n2309 & n18888;
  assign n18890 = ~n2306 & n18889;
  assign n18891 = ~n500 & n18890;
  assign n18892 = n2316 & n18891;
  assign n18893 = n3555 & n18892;
  assign n18894 = n3801 & n18893;
  assign n18895 = n3495 & n18894;
  assign n18896 = n3226 & n18895;
  assign n18897 = ~n3107 & n18896;
  assign n18898 = ~n3097 & n18897;
  assign n18899 = ~n3067 & n18898;
  assign n18900 = ~n3828 & n18565;
  assign n18901 = n3833 & n18900;
  assign n18902 = pi097 & ~n501;
  assign n18903 = n2311 & n18902;
  assign n18904 = n3813 & n18903;
  assign n18905 = n3811 & n18904;
  assign n18906 = ~n2306 & n18905;
  assign n18907 = n3819 & n18906;
  assign n18908 = n3823 & n18907;
  assign n18909 = n3809 & n18908;
  assign n18910 = ~n18901 & ~n18909;
  assign n18911 = ~n18899 & n18910;
  assign n18912 = pi073 & ~n2363;
  assign n18913 = n3847 & n18912;
  assign n18914 = n3855 & n18913;
  assign n18915 = n3843 & n18914;
  assign n18916 = n3869 & n18915;
  assign n18917 = ~n3066 & n18916;
  assign n18918 = n3874 & n18917;
  assign n18919 = ~n3837 & n18918;
  assign n18920 = n3903 & n18551;
  assign n18921 = n3907 & n18920;
  assign n18922 = ~n1372 & n18921;
  assign n18923 = ~n2243 & n18922;
  assign n18924 = ~n3104 & n18923;
  assign n18925 = ~n3901 & n18924;
  assign n18926 = ~n3837 & n18925;
  assign n18927 = ~n3900 & n18926;
  assign n18928 = ~n18919 & ~n18927;
  assign n18929 = pi081 & ~n3864;
  assign n18930 = ~n3919 & n18929;
  assign n18931 = ~n3916 & n18930;
  assign n18932 = n3924 & n18931;
  assign n18933 = ~n1897 & n18541;
  assign n18934 = n3082 & n18933;
  assign n18935 = n3888 & n18934;
  assign n18936 = ~n3886 & n18935;
  assign n18937 = n3885 & n18936;
  assign n18938 = ~n2242 & n18937;
  assign n18939 = ~n3095 & n18938;
  assign n18940 = ~n3878 & n18939;
  assign n18941 = ~n3877 & n18940;
  assign n18942 = ~n3837 & n18941;
  assign n18943 = ~n18932 & ~n18942;
  assign n18944 = n18928 & n18943;
  assign po050 = ~n18911 | ~n18944;
  assign n18946 = pi090 & ~n501;
  assign n18947 = n2311 & n18946;
  assign n18948 = n2309 & n18947;
  assign n18949 = ~n2306 & n18948;
  assign n18950 = ~n500 & n18949;
  assign n18951 = n2316 & n18950;
  assign n18952 = n3555 & n18951;
  assign n18953 = n3801 & n18952;
  assign n18954 = n3495 & n18953;
  assign n18955 = n3226 & n18954;
  assign n18956 = ~n3107 & n18955;
  assign n18957 = ~n3097 & n18956;
  assign n18958 = ~n3067 & n18957;
  assign n18959 = ~n3828 & n18603;
  assign n18960 = n3833 & n18959;
  assign n18961 = pi098 & ~n501;
  assign n18962 = n2311 & n18961;
  assign n18963 = n3813 & n18962;
  assign n18964 = n3811 & n18963;
  assign n18965 = ~n2306 & n18964;
  assign n18966 = n3819 & n18965;
  assign n18967 = n3823 & n18966;
  assign n18968 = n3809 & n18967;
  assign n18969 = ~n18960 & ~n18968;
  assign n18970 = ~n18958 & n18969;
  assign n18971 = pi074 & ~n2363;
  assign n18972 = n3847 & n18971;
  assign n18973 = n3855 & n18972;
  assign n18974 = n3843 & n18973;
  assign n18975 = n3869 & n18974;
  assign n18976 = ~n3066 & n18975;
  assign n18977 = n3874 & n18976;
  assign n18978 = ~n3837 & n18977;
  assign n18979 = n3903 & n18589;
  assign n18980 = n3907 & n18979;
  assign n18981 = ~n1372 & n18980;
  assign n18982 = ~n2243 & n18981;
  assign n18983 = ~n3104 & n18982;
  assign n18984 = ~n3901 & n18983;
  assign n18985 = ~n3837 & n18984;
  assign n18986 = ~n3900 & n18985;
  assign n18987 = ~n18978 & ~n18986;
  assign n18988 = pi082 & ~n3864;
  assign n18989 = ~n3919 & n18988;
  assign n18990 = ~n3916 & n18989;
  assign n18991 = n3924 & n18990;
  assign n18992 = ~n1897 & n18579;
  assign n18993 = n3082 & n18992;
  assign n18994 = n3888 & n18993;
  assign n18995 = ~n3886 & n18994;
  assign n18996 = n3885 & n18995;
  assign n18997 = ~n2242 & n18996;
  assign n18998 = ~n3095 & n18997;
  assign n18999 = ~n3878 & n18998;
  assign n19000 = ~n3877 & n18999;
  assign n19001 = ~n3837 & n19000;
  assign n19002 = ~n18991 & ~n19001;
  assign n19003 = n18987 & n19002;
  assign po051 = ~n18970 | ~n19003;
  assign n19005 = pi091 & ~n501;
  assign n19006 = n2311 & n19005;
  assign n19007 = n2309 & n19006;
  assign n19008 = ~n2306 & n19007;
  assign n19009 = ~n500 & n19008;
  assign n19010 = n2316 & n19009;
  assign n19011 = n3555 & n19010;
  assign n19012 = n3801 & n19011;
  assign n19013 = n3495 & n19012;
  assign n19014 = n3226 & n19013;
  assign n19015 = ~n3107 & n19014;
  assign n19016 = ~n3097 & n19015;
  assign n19017 = ~n3067 & n19016;
  assign n19018 = ~n3828 & n18641;
  assign n19019 = n3833 & n19018;
  assign n19020 = pi099 & ~n501;
  assign n19021 = n2311 & n19020;
  assign n19022 = n3813 & n19021;
  assign n19023 = n3811 & n19022;
  assign n19024 = ~n2306 & n19023;
  assign n19025 = n3819 & n19024;
  assign n19026 = n3823 & n19025;
  assign n19027 = n3809 & n19026;
  assign n19028 = ~n19019 & ~n19027;
  assign n19029 = ~n19017 & n19028;
  assign n19030 = pi075 & ~n2363;
  assign n19031 = n3847 & n19030;
  assign n19032 = n3855 & n19031;
  assign n19033 = n3843 & n19032;
  assign n19034 = n3869 & n19033;
  assign n19035 = ~n3066 & n19034;
  assign n19036 = n3874 & n19035;
  assign n19037 = ~n3837 & n19036;
  assign n19038 = n3903 & n18627;
  assign n19039 = n3907 & n19038;
  assign n19040 = ~n1372 & n19039;
  assign n19041 = ~n2243 & n19040;
  assign n19042 = ~n3104 & n19041;
  assign n19043 = ~n3901 & n19042;
  assign n19044 = ~n3837 & n19043;
  assign n19045 = ~n3900 & n19044;
  assign n19046 = ~n19037 & ~n19045;
  assign n19047 = pi083 & ~n3864;
  assign n19048 = ~n3919 & n19047;
  assign n19049 = ~n3916 & n19048;
  assign n19050 = n3924 & n19049;
  assign n19051 = ~n1897 & n18617;
  assign n19052 = n3082 & n19051;
  assign n19053 = n3888 & n19052;
  assign n19054 = ~n3886 & n19053;
  assign n19055 = n3885 & n19054;
  assign n19056 = ~n2242 & n19055;
  assign n19057 = ~n3095 & n19056;
  assign n19058 = ~n3878 & n19057;
  assign n19059 = ~n3877 & n19058;
  assign n19060 = ~n3837 & n19059;
  assign n19061 = ~n19050 & ~n19060;
  assign n19062 = n19046 & n19061;
  assign po052 = ~n19029 | ~n19062;
  assign n19064 = pi092 & ~n501;
  assign n19065 = n2311 & n19064;
  assign n19066 = n2309 & n19065;
  assign n19067 = ~n2306 & n19066;
  assign n19068 = ~n500 & n19067;
  assign n19069 = n2316 & n19068;
  assign n19070 = n3555 & n19069;
  assign n19071 = n3801 & n19070;
  assign n19072 = n3495 & n19071;
  assign n19073 = n3226 & n19072;
  assign n19074 = ~n3107 & n19073;
  assign n19075 = ~n3097 & n19074;
  assign n19076 = ~n3067 & n19075;
  assign n19077 = ~n3828 & n18679;
  assign n19078 = n3833 & n19077;
  assign n19079 = pi100 & ~n501;
  assign n19080 = n2311 & n19079;
  assign n19081 = n3813 & n19080;
  assign n19082 = n3811 & n19081;
  assign n19083 = ~n2306 & n19082;
  assign n19084 = n3819 & n19083;
  assign n19085 = n3823 & n19084;
  assign n19086 = n3809 & n19085;
  assign n19087 = ~n19078 & ~n19086;
  assign n19088 = ~n19076 & n19087;
  assign n19089 = pi076 & ~n2363;
  assign n19090 = n3847 & n19089;
  assign n19091 = n3855 & n19090;
  assign n19092 = n3843 & n19091;
  assign n19093 = n3869 & n19092;
  assign n19094 = ~n3066 & n19093;
  assign n19095 = n3874 & n19094;
  assign n19096 = ~n3837 & n19095;
  assign n19097 = n3903 & n18665;
  assign n19098 = n3907 & n19097;
  assign n19099 = ~n1372 & n19098;
  assign n19100 = ~n2243 & n19099;
  assign n19101 = ~n3104 & n19100;
  assign n19102 = ~n3901 & n19101;
  assign n19103 = ~n3837 & n19102;
  assign n19104 = ~n3900 & n19103;
  assign n19105 = ~n19096 & ~n19104;
  assign n19106 = pi084 & ~n3864;
  assign n19107 = ~n3919 & n19106;
  assign n19108 = ~n3916 & n19107;
  assign n19109 = n3924 & n19108;
  assign n19110 = ~n1897 & n18655;
  assign n19111 = n3082 & n19110;
  assign n19112 = n3888 & n19111;
  assign n19113 = ~n3886 & n19112;
  assign n19114 = n3885 & n19113;
  assign n19115 = ~n2242 & n19114;
  assign n19116 = ~n3095 & n19115;
  assign n19117 = ~n3878 & n19116;
  assign n19118 = ~n3877 & n19117;
  assign n19119 = ~n3837 & n19118;
  assign n19120 = ~n19109 & ~n19119;
  assign n19121 = n19105 & n19120;
  assign po053 = ~n19088 | ~n19121;
  assign n19123 = pi093 & ~n501;
  assign n19124 = n2311 & n19123;
  assign n19125 = n2309 & n19124;
  assign n19126 = ~n2306 & n19125;
  assign n19127 = ~n500 & n19126;
  assign n19128 = n2316 & n19127;
  assign n19129 = n3555 & n19128;
  assign n19130 = n3801 & n19129;
  assign n19131 = n3495 & n19130;
  assign n19132 = n3226 & n19131;
  assign n19133 = ~n3107 & n19132;
  assign n19134 = ~n3097 & n19133;
  assign n19135 = ~n3067 & n19134;
  assign n19136 = ~n3828 & n18717;
  assign n19137 = n3833 & n19136;
  assign n19138 = pi101 & ~n501;
  assign n19139 = n2311 & n19138;
  assign n19140 = n3813 & n19139;
  assign n19141 = n3811 & n19140;
  assign n19142 = ~n2306 & n19141;
  assign n19143 = n3819 & n19142;
  assign n19144 = n3823 & n19143;
  assign n19145 = n3809 & n19144;
  assign n19146 = ~n19137 & ~n19145;
  assign n19147 = ~n19135 & n19146;
  assign n19148 = pi077 & ~n2363;
  assign n19149 = n3847 & n19148;
  assign n19150 = n3855 & n19149;
  assign n19151 = n3843 & n19150;
  assign n19152 = n3869 & n19151;
  assign n19153 = ~n3066 & n19152;
  assign n19154 = n3874 & n19153;
  assign n19155 = ~n3837 & n19154;
  assign n19156 = n3903 & n18703;
  assign n19157 = n3907 & n19156;
  assign n19158 = ~n1372 & n19157;
  assign n19159 = ~n2243 & n19158;
  assign n19160 = ~n3104 & n19159;
  assign n19161 = ~n3901 & n19160;
  assign n19162 = ~n3837 & n19161;
  assign n19163 = ~n3900 & n19162;
  assign n19164 = ~n19155 & ~n19163;
  assign n19165 = pi085 & ~n3864;
  assign n19166 = ~n3919 & n19165;
  assign n19167 = ~n3916 & n19166;
  assign n19168 = n3924 & n19167;
  assign n19169 = ~n1897 & n18693;
  assign n19170 = n3082 & n19169;
  assign n19171 = n3888 & n19170;
  assign n19172 = ~n3886 & n19171;
  assign n19173 = n3885 & n19172;
  assign n19174 = ~n2242 & n19173;
  assign n19175 = ~n3095 & n19174;
  assign n19176 = ~n3878 & n19175;
  assign n19177 = ~n3877 & n19176;
  assign n19178 = ~n3837 & n19177;
  assign n19179 = ~n19168 & ~n19178;
  assign n19180 = n19164 & n19179;
  assign po054 = ~n19147 | ~n19180;
  assign n19182 = pi094 & ~n501;
  assign n19183 = n2311 & n19182;
  assign n19184 = n2309 & n19183;
  assign n19185 = ~n2306 & n19184;
  assign n19186 = ~n500 & n19185;
  assign n19187 = n2316 & n19186;
  assign n19188 = n3555 & n19187;
  assign n19189 = n3801 & n19188;
  assign n19190 = n3495 & n19189;
  assign n19191 = n3226 & n19190;
  assign n19192 = ~n3107 & n19191;
  assign n19193 = ~n3097 & n19192;
  assign n19194 = ~n3067 & n19193;
  assign n19195 = ~n3828 & n18755;
  assign n19196 = n3833 & n19195;
  assign n19197 = pi102 & ~n501;
  assign n19198 = n2311 & n19197;
  assign n19199 = n3813 & n19198;
  assign n19200 = n3811 & n19199;
  assign n19201 = ~n2306 & n19200;
  assign n19202 = n3819 & n19201;
  assign n19203 = n3823 & n19202;
  assign n19204 = n3809 & n19203;
  assign n19205 = ~n19196 & ~n19204;
  assign n19206 = ~n19194 & n19205;
  assign n19207 = pi078 & ~n2363;
  assign n19208 = n3847 & n19207;
  assign n19209 = n3855 & n19208;
  assign n19210 = n3843 & n19209;
  assign n19211 = n3869 & n19210;
  assign n19212 = ~n3066 & n19211;
  assign n19213 = n3874 & n19212;
  assign n19214 = ~n3837 & n19213;
  assign n19215 = n3903 & n18741;
  assign n19216 = n3907 & n19215;
  assign n19217 = ~n1372 & n19216;
  assign n19218 = ~n2243 & n19217;
  assign n19219 = ~n3104 & n19218;
  assign n19220 = ~n3901 & n19219;
  assign n19221 = ~n3837 & n19220;
  assign n19222 = ~n3900 & n19221;
  assign n19223 = ~n19214 & ~n19222;
  assign n19224 = pi086 & ~n3864;
  assign n19225 = ~n3919 & n19224;
  assign n19226 = ~n3916 & n19225;
  assign n19227 = n3924 & n19226;
  assign n19228 = ~n1897 & n18731;
  assign n19229 = n3082 & n19228;
  assign n19230 = n3888 & n19229;
  assign n19231 = ~n3886 & n19230;
  assign n19232 = n3885 & n19231;
  assign n19233 = ~n2242 & n19232;
  assign n19234 = ~n3095 & n19233;
  assign n19235 = ~n3878 & n19234;
  assign n19236 = ~n3877 & n19235;
  assign n19237 = ~n3837 & n19236;
  assign n19238 = ~n19227 & ~n19237;
  assign n19239 = n19223 & n19238;
  assign po055 = ~n19206 | ~n19239;
  assign n19241 = n2633 & n18794;
  assign n19242 = n3977 & n19241;
  assign n19243 = n4074 & n19242;
  assign n19244 = n2936 & n19243;
  assign n19245 = ~n4004 & n19244;
  assign n19246 = ~n3066 & n19245;
  assign n19247 = ~n3983 & n19246;
  assign n19248 = ~n4003 & n19247;
  assign n19249 = n4023 & n19248;
  assign n19250 = n3883 & n5837;
  assign n19251 = n3882 & n19250;
  assign n19252 = pi055 & ~n2077;
  assign n19253 = ~n2078 & n19252;
  assign n19254 = ~n2076 & n19253;
  assign n19255 = ~n2143 & n19254;
  assign n19256 = n2207 & n19255;
  assign n19257 = n1928 & n19256;
  assign n19258 = n4827 & n19257;
  assign n19259 = n19251 & n19258;
  assign n19260 = ~n4025 & n19259;
  assign n19261 = ~n2242 & n19260;
  assign n19262 = ~n3095 & n19261;
  assign n19263 = ~n3997 & n19262;
  assign n19264 = ~n4003 & n19263;
  assign n19265 = n4044 & n19264;
  assign n19266 = ~n19249 & ~n19265;
  assign n19267 = pi039 & ~n1169;
  assign n19268 = ~n1170 & n19267;
  assign n19269 = ~n1168 & n19268;
  assign n19270 = ~n1144 & n19269;
  assign n19271 = ~n1115 & n19270;
  assign n19272 = ~n1086 & n19271;
  assign n19273 = n1057 & n19272;
  assign n19274 = n1239 & n19273;
  assign n19275 = n843 & n19274;
  assign n19276 = n720 & n19275;
  assign n19277 = n4048 & n19276;
  assign n19278 = ~n4047 & n19277;
  assign n19279 = n3831 & n19278;
  assign n19280 = ~n3104 & n19279;
  assign n19281 = ~n3971 & n19280;
  assign n19282 = ~n4003 & n19281;
  assign n19283 = n4871 & n19282;
  assign n19284 = ~n3931 & n18813;
  assign n19285 = ~n4070 & n19284;
  assign n19286 = ~n4068 & n19285;
  assign n19287 = n4842 & n19286;
  assign n19288 = ~n19283 & ~n19287;
  assign n19289 = n19266 & n19288;
  assign n19290 = pi095 & ~po149;
  assign n19291 = ~n3932 & n19290;
  assign n19292 = n4127 & n19291;
  assign n19293 = pi111 & ~n501;
  assign n19294 = n4792 & n19293;
  assign n19295 = n4790 & n19294;
  assign n19296 = n4800 & n19295;
  assign n19297 = ~n996 & n19296;
  assign n19298 = ~n2306 & n19297;
  assign n19299 = n3819 & n19298;
  assign n19300 = n4789 & n19299;
  assign n19301 = n3823 & n19300;
  assign n19302 = n4787 & n19301;
  assign n19303 = ~n19292 & ~n19302;
  assign n19304 = pi103 & ~n501;
  assign n19305 = n2311 & n19304;
  assign n19306 = n3813 & n19305;
  assign n19307 = n3811 & n19306;
  assign n19308 = ~n2306 & n19307;
  assign n19309 = n3819 & n19308;
  assign n19310 = n3823 & n19309;
  assign n19311 = n4770 & n19310;
  assign n19312 = n4612 & n19311;
  assign n19313 = n4253 & n19312;
  assign n19314 = ~n4134 & n19313;
  assign n19315 = n4784 & n19314;
  assign n19316 = pi087 & ~n3251;
  assign n19317 = ~n3252 & n19316;
  assign n19318 = ~n3250 & n19317;
  assign n19319 = ~n3524 & n19318;
  assign n19320 = n4095 & n19319;
  assign n19321 = n5062 & n19320;
  assign n19322 = n5068 & n19321;
  assign n19323 = n3226 & n19322;
  assign n19324 = ~n3950 & n19323;
  assign n19325 = ~n3940 & n19324;
  assign n19326 = ~n3932 & n19325;
  assign n19327 = n4000 & n19326;
  assign n19328 = ~n19315 & ~n19327;
  assign n19329 = n19303 & n19328;
  assign po056 = ~n19289 | ~n19329;
  assign n19331 = n4030 & n18862;
  assign n19332 = n4029 & n19331;
  assign n19333 = ~n4025 & n19332;
  assign n19334 = ~n2242 & n19333;
  assign n19335 = ~n3095 & n19334;
  assign n19336 = ~n3997 & n19335;
  assign n19337 = ~n4003 & n19336;
  assign n19338 = n4044 & n19337;
  assign n19339 = pi104 & ~n501;
  assign n19340 = n2311 & n19339;
  assign n19341 = n3813 & n19340;
  assign n19342 = n3811 & n19341;
  assign n19343 = ~n2306 & n19342;
  assign n19344 = n3819 & n19343;
  assign n19345 = n3823 & n19344;
  assign n19346 = n4770 & n19345;
  assign n19347 = n4612 & n19346;
  assign n19348 = n4253 & n19347;
  assign n19349 = ~n4134 & n19348;
  assign n19350 = n4784 & n19349;
  assign n19351 = ~n19338 & ~n19350;
  assign n19352 = pi096 & ~po149;
  assign n19353 = ~n3932 & n19352;
  assign n19354 = n4127 & n19353;
  assign n19355 = n2633 & n18828;
  assign n19356 = n3977 & n19355;
  assign n19357 = n4074 & n19356;
  assign n19358 = n2936 & n19357;
  assign n19359 = ~n4004 & n19358;
  assign n19360 = ~n3066 & n19359;
  assign n19361 = ~n3983 & n19360;
  assign n19362 = ~n4003 & n19361;
  assign n19363 = n4023 & n19362;
  assign n19364 = ~n19354 & ~n19363;
  assign n19365 = n19351 & n19364;
  assign n19366 = n843 & n18172;
  assign n19367 = n720 & n19366;
  assign n19368 = n4048 & n19367;
  assign n19369 = ~n4047 & n19368;
  assign n19370 = n3831 & n19369;
  assign n19371 = ~n3104 & n19370;
  assign n19372 = ~n3971 & n19371;
  assign n19373 = ~n4003 & n19372;
  assign n19374 = n4871 & n19373;
  assign n19375 = pi112 & ~n501;
  assign n19376 = n4792 & n19375;
  assign n19377 = n4790 & n19376;
  assign n19378 = n4800 & n19377;
  assign n19379 = ~n996 & n19378;
  assign n19380 = ~n2306 & n19379;
  assign n19381 = n3819 & n19380;
  assign n19382 = n4789 & n19381;
  assign n19383 = n3823 & n19382;
  assign n19384 = n4787 & n19383;
  assign n19385 = ~n19374 & ~n19384;
  assign n19386 = pi088 & ~n3524;
  assign n19387 = n4097 & n19386;
  assign n19388 = n4105 & n19387;
  assign n19389 = n4093 & n19388;
  assign n19390 = n4088 & n19389;
  assign n19391 = ~n3950 & n19390;
  assign n19392 = ~n3940 & n19391;
  assign n19393 = ~n3932 & n19392;
  assign n19394 = n4000 & n19393;
  assign n19395 = ~n3931 & n18880;
  assign n19396 = ~n4070 & n19395;
  assign n19397 = ~n4068 & n19396;
  assign n19398 = n4842 & n19397;
  assign n19399 = ~n19394 & ~n19398;
  assign n19400 = n19385 & n19399;
  assign po057 = ~n19365 | ~n19400;
  assign n19402 = n4030 & n18934;
  assign n19403 = n4029 & n19402;
  assign n19404 = ~n4025 & n19403;
  assign n19405 = ~n2242 & n19404;
  assign n19406 = ~n3095 & n19405;
  assign n19407 = ~n3997 & n19406;
  assign n19408 = ~n4003 & n19407;
  assign n19409 = n4044 & n19408;
  assign n19410 = pi105 & ~n501;
  assign n19411 = n2311 & n19410;
  assign n19412 = n3813 & n19411;
  assign n19413 = n3811 & n19412;
  assign n19414 = ~n2306 & n19413;
  assign n19415 = n3819 & n19414;
  assign n19416 = n3823 & n19415;
  assign n19417 = n4770 & n19416;
  assign n19418 = n4612 & n19417;
  assign n19419 = n4253 & n19418;
  assign n19420 = ~n4134 & n19419;
  assign n19421 = n4784 & n19420;
  assign n19422 = ~n19409 & ~n19421;
  assign n19423 = pi097 & ~po149;
  assign n19424 = ~n3932 & n19423;
  assign n19425 = n4127 & n19424;
  assign n19426 = n2633 & n18912;
  assign n19427 = n3977 & n19426;
  assign n19428 = n4074 & n19427;
  assign n19429 = n2936 & n19428;
  assign n19430 = ~n4004 & n19429;
  assign n19431 = ~n3066 & n19430;
  assign n19432 = ~n3983 & n19431;
  assign n19433 = ~n4003 & n19432;
  assign n19434 = n4023 & n19433;
  assign n19435 = ~n19425 & ~n19434;
  assign n19436 = n19422 & n19435;
  assign n19437 = pi089 & ~n3524;
  assign n19438 = n4097 & n19437;
  assign n19439 = n4105 & n19438;
  assign n19440 = n4093 & n19439;
  assign n19441 = n4088 & n19440;
  assign n19442 = ~n3950 & n19441;
  assign n19443 = ~n3940 & n19442;
  assign n19444 = ~n3932 & n19443;
  assign n19445 = n4000 & n19444;
  assign n19446 = pi113 & ~n501;
  assign n19447 = n4792 & n19446;
  assign n19448 = n4790 & n19447;
  assign n19449 = n4800 & n19448;
  assign n19450 = ~n996 & n19449;
  assign n19451 = ~n2306 & n19450;
  assign n19452 = n3819 & n19451;
  assign n19453 = n4789 & n19452;
  assign n19454 = n3823 & n19453;
  assign n19455 = n4787 & n19454;
  assign n19456 = ~n19445 & ~n19455;
  assign n19457 = n843 & n18184;
  assign n19458 = n720 & n19457;
  assign n19459 = n4048 & n19458;
  assign n19460 = ~n4047 & n19459;
  assign n19461 = n3831 & n19460;
  assign n19462 = ~n3104 & n19461;
  assign n19463 = ~n3971 & n19462;
  assign n19464 = ~n4003 & n19463;
  assign n19465 = n4871 & n19464;
  assign n19466 = ~n3931 & n18929;
  assign n19467 = ~n4070 & n19466;
  assign n19468 = ~n4068 & n19467;
  assign n19469 = n4842 & n19468;
  assign n19470 = ~n19465 & ~n19469;
  assign n19471 = n19456 & n19470;
  assign po058 = ~n19436 | ~n19471;
  assign n19473 = n4030 & n18993;
  assign n19474 = n4029 & n19473;
  assign n19475 = ~n4025 & n19474;
  assign n19476 = ~n2242 & n19475;
  assign n19477 = ~n3095 & n19476;
  assign n19478 = ~n3997 & n19477;
  assign n19479 = ~n4003 & n19478;
  assign n19480 = n4044 & n19479;
  assign n19481 = pi106 & ~n501;
  assign n19482 = n2311 & n19481;
  assign n19483 = n3813 & n19482;
  assign n19484 = n3811 & n19483;
  assign n19485 = ~n2306 & n19484;
  assign n19486 = n3819 & n19485;
  assign n19487 = n3823 & n19486;
  assign n19488 = n4770 & n19487;
  assign n19489 = n4612 & n19488;
  assign n19490 = n4253 & n19489;
  assign n19491 = ~n4134 & n19490;
  assign n19492 = n4784 & n19491;
  assign n19493 = ~n19480 & ~n19492;
  assign n19494 = pi098 & ~po149;
  assign n19495 = ~n3932 & n19494;
  assign n19496 = n4127 & n19495;
  assign n19497 = n2633 & n18971;
  assign n19498 = n3977 & n19497;
  assign n19499 = n4074 & n19498;
  assign n19500 = n2936 & n19499;
  assign n19501 = ~n4004 & n19500;
  assign n19502 = ~n3066 & n19501;
  assign n19503 = ~n3983 & n19502;
  assign n19504 = ~n4003 & n19503;
  assign n19505 = n4023 & n19504;
  assign n19506 = ~n19496 & ~n19505;
  assign n19507 = n19493 & n19506;
  assign n19508 = pi090 & ~n3524;
  assign n19509 = n4097 & n19508;
  assign n19510 = n4105 & n19509;
  assign n19511 = n4093 & n19510;
  assign n19512 = n4088 & n19511;
  assign n19513 = ~n3950 & n19512;
  assign n19514 = ~n3940 & n19513;
  assign n19515 = ~n3932 & n19514;
  assign n19516 = n4000 & n19515;
  assign n19517 = pi114 & ~n501;
  assign n19518 = n4792 & n19517;
  assign n19519 = n4790 & n19518;
  assign n19520 = n4800 & n19519;
  assign n19521 = ~n996 & n19520;
  assign n19522 = ~n2306 & n19521;
  assign n19523 = n3819 & n19522;
  assign n19524 = n4789 & n19523;
  assign n19525 = n3823 & n19524;
  assign n19526 = n4787 & n19525;
  assign n19527 = ~n19516 & ~n19526;
  assign n19528 = n843 & n18196;
  assign n19529 = n720 & n19528;
  assign n19530 = n4048 & n19529;
  assign n19531 = ~n4047 & n19530;
  assign n19532 = n3831 & n19531;
  assign n19533 = ~n3104 & n19532;
  assign n19534 = ~n3971 & n19533;
  assign n19535 = ~n4003 & n19534;
  assign n19536 = n4871 & n19535;
  assign n19537 = ~n3931 & n18988;
  assign n19538 = ~n4070 & n19537;
  assign n19539 = ~n4068 & n19538;
  assign n19540 = n4842 & n19539;
  assign n19541 = ~n19536 & ~n19540;
  assign n19542 = n19527 & n19541;
  assign po059 = ~n19507 | ~n19542;
  assign n19544 = n4030 & n19052;
  assign n19545 = n4029 & n19544;
  assign n19546 = ~n4025 & n19545;
  assign n19547 = ~n2242 & n19546;
  assign n19548 = ~n3095 & n19547;
  assign n19549 = ~n3997 & n19548;
  assign n19550 = ~n4003 & n19549;
  assign n19551 = n4044 & n19550;
  assign n19552 = pi107 & ~n501;
  assign n19553 = n2311 & n19552;
  assign n19554 = n3813 & n19553;
  assign n19555 = n3811 & n19554;
  assign n19556 = ~n2306 & n19555;
  assign n19557 = n3819 & n19556;
  assign n19558 = n3823 & n19557;
  assign n19559 = n4770 & n19558;
  assign n19560 = n4612 & n19559;
  assign n19561 = n4253 & n19560;
  assign n19562 = ~n4134 & n19561;
  assign n19563 = n4784 & n19562;
  assign n19564 = ~n19551 & ~n19563;
  assign n19565 = pi099 & ~po149;
  assign n19566 = ~n3932 & n19565;
  assign n19567 = n4127 & n19566;
  assign n19568 = n2633 & n19030;
  assign n19569 = n3977 & n19568;
  assign n19570 = n4074 & n19569;
  assign n19571 = n2936 & n19570;
  assign n19572 = ~n4004 & n19571;
  assign n19573 = ~n3066 & n19572;
  assign n19574 = ~n3983 & n19573;
  assign n19575 = ~n4003 & n19574;
  assign n19576 = n4023 & n19575;
  assign n19577 = ~n19567 & ~n19576;
  assign n19578 = n19564 & n19577;
  assign n19579 = pi091 & ~n3524;
  assign n19580 = n4097 & n19579;
  assign n19581 = n4105 & n19580;
  assign n19582 = n4093 & n19581;
  assign n19583 = n4088 & n19582;
  assign n19584 = ~n3950 & n19583;
  assign n19585 = ~n3940 & n19584;
  assign n19586 = ~n3932 & n19585;
  assign n19587 = n4000 & n19586;
  assign n19588 = pi115 & ~n501;
  assign n19589 = n4792 & n19588;
  assign n19590 = n4790 & n19589;
  assign n19591 = n4800 & n19590;
  assign n19592 = ~n996 & n19591;
  assign n19593 = ~n2306 & n19592;
  assign n19594 = n3819 & n19593;
  assign n19595 = n4789 & n19594;
  assign n19596 = n3823 & n19595;
  assign n19597 = n4787 & n19596;
  assign n19598 = ~n19587 & ~n19597;
  assign n19599 = n843 & n18208;
  assign n19600 = n720 & n19599;
  assign n19601 = n4048 & n19600;
  assign n19602 = ~n4047 & n19601;
  assign n19603 = n3831 & n19602;
  assign n19604 = ~n3104 & n19603;
  assign n19605 = ~n3971 & n19604;
  assign n19606 = ~n4003 & n19605;
  assign n19607 = n4871 & n19606;
  assign n19608 = ~n3931 & n19047;
  assign n19609 = ~n4070 & n19608;
  assign n19610 = ~n4068 & n19609;
  assign n19611 = n4842 & n19610;
  assign n19612 = ~n19607 & ~n19611;
  assign n19613 = n19598 & n19612;
  assign po060 = ~n19578 | ~n19613;
  assign n19615 = n4030 & n19111;
  assign n19616 = n4029 & n19615;
  assign n19617 = ~n4025 & n19616;
  assign n19618 = ~n2242 & n19617;
  assign n19619 = ~n3095 & n19618;
  assign n19620 = ~n3997 & n19619;
  assign n19621 = ~n4003 & n19620;
  assign n19622 = n4044 & n19621;
  assign n19623 = pi108 & ~n501;
  assign n19624 = n2311 & n19623;
  assign n19625 = n3813 & n19624;
  assign n19626 = n3811 & n19625;
  assign n19627 = ~n2306 & n19626;
  assign n19628 = n3819 & n19627;
  assign n19629 = n3823 & n19628;
  assign n19630 = n4770 & n19629;
  assign n19631 = n4612 & n19630;
  assign n19632 = n4253 & n19631;
  assign n19633 = ~n4134 & n19632;
  assign n19634 = n4784 & n19633;
  assign n19635 = ~n19622 & ~n19634;
  assign n19636 = pi100 & ~po149;
  assign n19637 = ~n3932 & n19636;
  assign n19638 = n4127 & n19637;
  assign n19639 = n2633 & n19089;
  assign n19640 = n3977 & n19639;
  assign n19641 = n4074 & n19640;
  assign n19642 = n2936 & n19641;
  assign n19643 = ~n4004 & n19642;
  assign n19644 = ~n3066 & n19643;
  assign n19645 = ~n3983 & n19644;
  assign n19646 = ~n4003 & n19645;
  assign n19647 = n4023 & n19646;
  assign n19648 = ~n19638 & ~n19647;
  assign n19649 = n19635 & n19648;
  assign n19650 = pi092 & ~n3524;
  assign n19651 = n4097 & n19650;
  assign n19652 = n4105 & n19651;
  assign n19653 = n4093 & n19652;
  assign n19654 = n4088 & n19653;
  assign n19655 = ~n3950 & n19654;
  assign n19656 = ~n3940 & n19655;
  assign n19657 = ~n3932 & n19656;
  assign n19658 = n4000 & n19657;
  assign n19659 = pi116 & ~n501;
  assign n19660 = n4792 & n19659;
  assign n19661 = n4790 & n19660;
  assign n19662 = n4800 & n19661;
  assign n19663 = ~n996 & n19662;
  assign n19664 = ~n2306 & n19663;
  assign n19665 = n3819 & n19664;
  assign n19666 = n4789 & n19665;
  assign n19667 = n3823 & n19666;
  assign n19668 = n4787 & n19667;
  assign n19669 = ~n19658 & ~n19668;
  assign n19670 = n843 & n18220;
  assign n19671 = n720 & n19670;
  assign n19672 = n4048 & n19671;
  assign n19673 = ~n4047 & n19672;
  assign n19674 = n3831 & n19673;
  assign n19675 = ~n3104 & n19674;
  assign n19676 = ~n3971 & n19675;
  assign n19677 = ~n4003 & n19676;
  assign n19678 = n4871 & n19677;
  assign n19679 = ~n3931 & n19106;
  assign n19680 = ~n4070 & n19679;
  assign n19681 = ~n4068 & n19680;
  assign n19682 = n4842 & n19681;
  assign n19683 = ~n19678 & ~n19682;
  assign n19684 = n19669 & n19683;
  assign po061 = ~n19649 | ~n19684;
  assign n19686 = n4030 & n19170;
  assign n19687 = n4029 & n19686;
  assign n19688 = ~n4025 & n19687;
  assign n19689 = ~n2242 & n19688;
  assign n19690 = ~n3095 & n19689;
  assign n19691 = ~n3997 & n19690;
  assign n19692 = ~n4003 & n19691;
  assign n19693 = n4044 & n19692;
  assign n19694 = pi109 & ~n501;
  assign n19695 = n2311 & n19694;
  assign n19696 = n3813 & n19695;
  assign n19697 = n3811 & n19696;
  assign n19698 = ~n2306 & n19697;
  assign n19699 = n3819 & n19698;
  assign n19700 = n3823 & n19699;
  assign n19701 = n4770 & n19700;
  assign n19702 = n4612 & n19701;
  assign n19703 = n4253 & n19702;
  assign n19704 = ~n4134 & n19703;
  assign n19705 = n4784 & n19704;
  assign n19706 = ~n19693 & ~n19705;
  assign n19707 = pi101 & ~po149;
  assign n19708 = ~n3932 & n19707;
  assign n19709 = n4127 & n19708;
  assign n19710 = n2633 & n19148;
  assign n19711 = n3977 & n19710;
  assign n19712 = n4074 & n19711;
  assign n19713 = n2936 & n19712;
  assign n19714 = ~n4004 & n19713;
  assign n19715 = ~n3066 & n19714;
  assign n19716 = ~n3983 & n19715;
  assign n19717 = ~n4003 & n19716;
  assign n19718 = n4023 & n19717;
  assign n19719 = ~n19709 & ~n19718;
  assign n19720 = n19706 & n19719;
  assign n19721 = pi093 & ~n3524;
  assign n19722 = n4097 & n19721;
  assign n19723 = n4105 & n19722;
  assign n19724 = n4093 & n19723;
  assign n19725 = n4088 & n19724;
  assign n19726 = ~n3950 & n19725;
  assign n19727 = ~n3940 & n19726;
  assign n19728 = ~n3932 & n19727;
  assign n19729 = n4000 & n19728;
  assign n19730 = pi117 & ~n501;
  assign n19731 = n4792 & n19730;
  assign n19732 = n4790 & n19731;
  assign n19733 = n4800 & n19732;
  assign n19734 = ~n996 & n19733;
  assign n19735 = ~n2306 & n19734;
  assign n19736 = n3819 & n19735;
  assign n19737 = n4789 & n19736;
  assign n19738 = n3823 & n19737;
  assign n19739 = n4787 & n19738;
  assign n19740 = ~n19729 & ~n19739;
  assign n19741 = n843 & n18232;
  assign n19742 = n720 & n19741;
  assign n19743 = n4048 & n19742;
  assign n19744 = ~n4047 & n19743;
  assign n19745 = n3831 & n19744;
  assign n19746 = ~n3104 & n19745;
  assign n19747 = ~n3971 & n19746;
  assign n19748 = ~n4003 & n19747;
  assign n19749 = n4871 & n19748;
  assign n19750 = ~n3931 & n19165;
  assign n19751 = ~n4070 & n19750;
  assign n19752 = ~n4068 & n19751;
  assign n19753 = n4842 & n19752;
  assign n19754 = ~n19749 & ~n19753;
  assign n19755 = n19740 & n19754;
  assign po062 = ~n19720 | ~n19755;
  assign n19757 = n4030 & n19229;
  assign n19758 = n4029 & n19757;
  assign n19759 = ~n4025 & n19758;
  assign n19760 = ~n2242 & n19759;
  assign n19761 = ~n3095 & n19760;
  assign n19762 = ~n3997 & n19761;
  assign n19763 = ~n4003 & n19762;
  assign n19764 = n4044 & n19763;
  assign n19765 = pi110 & ~n501;
  assign n19766 = n2311 & n19765;
  assign n19767 = n3813 & n19766;
  assign n19768 = n3811 & n19767;
  assign n19769 = ~n2306 & n19768;
  assign n19770 = n3819 & n19769;
  assign n19771 = n3823 & n19770;
  assign n19772 = n4770 & n19771;
  assign n19773 = n4612 & n19772;
  assign n19774 = n4253 & n19773;
  assign n19775 = ~n4134 & n19774;
  assign n19776 = n4784 & n19775;
  assign n19777 = ~n19764 & ~n19776;
  assign n19778 = pi102 & ~po149;
  assign n19779 = ~n3932 & n19778;
  assign n19780 = n4127 & n19779;
  assign n19781 = n2633 & n19207;
  assign n19782 = n3977 & n19781;
  assign n19783 = n4074 & n19782;
  assign n19784 = n2936 & n19783;
  assign n19785 = ~n4004 & n19784;
  assign n19786 = ~n3066 & n19785;
  assign n19787 = ~n3983 & n19786;
  assign n19788 = ~n4003 & n19787;
  assign n19789 = n4023 & n19788;
  assign n19790 = ~n19780 & ~n19789;
  assign n19791 = n19777 & n19790;
  assign n19792 = pi094 & ~n3524;
  assign n19793 = n4097 & n19792;
  assign n19794 = n4105 & n19793;
  assign n19795 = n4093 & n19794;
  assign n19796 = n4088 & n19795;
  assign n19797 = ~n3950 & n19796;
  assign n19798 = ~n3940 & n19797;
  assign n19799 = ~n3932 & n19798;
  assign n19800 = n4000 & n19799;
  assign n19801 = pi118 & ~n501;
  assign n19802 = n4792 & n19801;
  assign n19803 = n4790 & n19802;
  assign n19804 = n4800 & n19803;
  assign n19805 = ~n996 & n19804;
  assign n19806 = ~n2306 & n19805;
  assign n19807 = n3819 & n19806;
  assign n19808 = n4789 & n19807;
  assign n19809 = n3823 & n19808;
  assign n19810 = n4787 & n19809;
  assign n19811 = ~n19800 & ~n19810;
  assign n19812 = n843 & n18244;
  assign n19813 = n720 & n19812;
  assign n19814 = n4048 & n19813;
  assign n19815 = ~n4047 & n19814;
  assign n19816 = n3831 & n19815;
  assign n19817 = ~n3104 & n19816;
  assign n19818 = ~n3971 & n19817;
  assign n19819 = ~n4003 & n19818;
  assign n19820 = n4871 & n19819;
  assign n19821 = ~n3931 & n19224;
  assign n19822 = ~n4070 & n19821;
  assign n19823 = ~n4068 & n19822;
  assign n19824 = n4842 & n19823;
  assign n19825 = ~n19820 & ~n19824;
  assign n19826 = n19811 & n19825;
  assign po063 = ~n19791 | ~n19826;
  assign n19828 = pi119 & ~n501;
  assign n19829 = n4792 & n19828;
  assign n19830 = n4790 & n19829;
  assign n19831 = n4800 & n19830;
  assign n19832 = ~n996 & n19831;
  assign n19833 = ~n2306 & n19832;
  assign n19834 = n3819 & n19833;
  assign n19835 = n4789 & n19834;
  assign n19836 = n3823 & n19835;
  assign n19837 = n5689 & n19836;
  assign n19838 = n5560 & n19837;
  assign n19839 = n5201 & n19838;
  assign n19840 = ~n5112 & n19839;
  assign n19841 = n5710 & n19840;
  assign n19842 = n2573 & n18794;
  assign n19843 = n5002 & n19842;
  assign n19844 = n5010 & n19843;
  assign n19845 = n4983 & n19844;
  assign n19846 = ~n4981 & n19845;
  assign n19847 = ~n3066 & n19846;
  assign n19848 = ~n3983 & n19847;
  assign n19849 = ~n4003 & n19848;
  assign n19850 = ~n4024 & n19849;
  assign n19851 = ~n4980 & n19850;
  assign n19852 = n4997 & n19851;
  assign n19853 = n4979 & n19852;
  assign n19854 = n1056 & n19271;
  assign n19855 = ~n1208 & n19854;
  assign n19856 = n4920 & n19855;
  assign n19857 = n4925 & n19856;
  assign n19858 = n4932 & n19857;
  assign n19859 = ~n4917 & n19858;
  assign n19860 = ~n1372 & n19859;
  assign n19861 = ~n2243 & n19860;
  assign n19862 = ~n3104 & n19861;
  assign n19863 = ~n3971 & n19862;
  assign n19864 = ~n4003 & n19863;
  assign n19865 = ~n4872 & n19864;
  assign n19866 = ~n4916 & n19865;
  assign n19867 = n4944 & n19866;
  assign n19868 = n4915 & n19867;
  assign n19869 = ~n19853 & ~n19868;
  assign n19870 = ~n19841 & n19869;
  assign n19871 = n5810 & n19250;
  assign n19872 = n4959 & n19257;
  assign n19873 = n19871 & n19872;
  assign n19874 = ~n4953 & n19873;
  assign n19875 = ~n2242 & n19874;
  assign n19876 = ~n3095 & n19875;
  assign n19877 = ~n3997 & n19876;
  assign n19878 = ~n4003 & n19877;
  assign n19879 = ~n4837 & n19878;
  assign n19880 = ~n4952 & n19879;
  assign n19881 = n4972 & n19880;
  assign n19882 = n4951 & n19881;
  assign n19883 = ~n4003 & n19284;
  assign n19884 = ~n4844 & n19883;
  assign n19885 = ~n4903 & n19884;
  assign n19886 = n4909 & n19885;
  assign n19887 = pi127 & ~n501;
  assign n19888 = n5714 & n19887;
  assign n19889 = n5725 & n19888;
  assign n19890 = ~n1172 & n19889;
  assign n19891 = ~n996 & n19890;
  assign n19892 = ~n2306 & n19891;
  assign n19893 = n3819 & n19892;
  assign n19894 = n3821 & n19893;
  assign n19895 = n5736 & n19894;
  assign n19896 = ~n1493 & n14226;
  assign n19897 = n5740 & n19896;
  assign n19898 = n19895 & n19897;
  assign n19899 = ~n19886 & ~n19898;
  assign n19900 = ~n19882 & n19899;
  assign n19901 = pi103 & ~n4644;
  assign n19902 = ~n4645 & n19901;
  assign n19903 = ~n4643 & n19902;
  assign n19904 = ~n4677 & n19903;
  assign n19905 = n4737 & n19904;
  assign n19906 = n4491 & n19905;
  assign n19907 = n4893 & n19906;
  assign n19908 = n4889 & n19907;
  assign n19909 = ~n4887 & n19908;
  assign n19910 = ~n4817 & n19909;
  assign n19911 = ~n4845 & n19910;
  assign n19912 = n4900 & n19911;
  assign n19913 = n4886 & n19912;
  assign n19914 = pi087 & ~n3524;
  assign n19915 = n4095 & n19914;
  assign n19916 = n5062 & n19915;
  assign n19917 = n5068 & n19916;
  assign n19918 = n5029 & n19917;
  assign n19919 = ~n5028 & n19918;
  assign n19920 = ~n3940 & n19919;
  assign n19921 = ~n4001 & n19920;
  assign n19922 = ~n4845 & n19921;
  assign n19923 = n5041 & n19922;
  assign n19924 = n5027 & n19923;
  assign n19925 = ~n19913 & ~n19924;
  assign n19926 = pi111 & ~n4858;
  assign n19927 = ~n4845 & n19926;
  assign n19928 = ~n4841 & n19927;
  assign n19929 = n4879 & n19928;
  assign n19930 = n4823 & n19929;
  assign n19931 = ~n4128 & n19290;
  assign n19932 = ~n4845 & n19931;
  assign n19933 = n5057 & n19932;
  assign n19934 = ~n19930 & ~n19933;
  assign n19935 = n19925 & n19934;
  assign n19936 = n19900 & n19935;
  assign po064 = ~n19870 | ~n19936;
  assign n19938 = n2573 & n18828;
  assign n19939 = n5002 & n19938;
  assign n19940 = n5010 & n19939;
  assign n19941 = n4983 & n19940;
  assign n19942 = ~n4981 & n19941;
  assign n19943 = ~n3066 & n19942;
  assign n19944 = ~n3983 & n19943;
  assign n19945 = ~n4003 & n19944;
  assign n19946 = ~n4024 & n19945;
  assign n19947 = ~n4980 & n19946;
  assign n19948 = n4997 & n19947;
  assign n19949 = n4979 & n19948;
  assign n19950 = n1928 & n18504;
  assign n19951 = n4959 & n19950;
  assign n19952 = n4958 & n19951;
  assign n19953 = ~n4953 & n19952;
  assign n19954 = ~n2242 & n19953;
  assign n19955 = ~n3095 & n19954;
  assign n19956 = ~n3997 & n19955;
  assign n19957 = ~n4003 & n19956;
  assign n19958 = ~n4837 & n19957;
  assign n19959 = ~n4952 & n19958;
  assign n19960 = n4972 & n19959;
  assign n19961 = n4951 & n19960;
  assign n19962 = pi104 & ~n4648;
  assign n19963 = n5087 & n19962;
  assign n19964 = n5085 & n19963;
  assign n19965 = n5097 & n19964;
  assign n19966 = n4889 & n19965;
  assign n19967 = ~n4887 & n19966;
  assign n19968 = ~n4817 & n19967;
  assign n19969 = ~n4845 & n19968;
  assign n19970 = n4900 & n19969;
  assign n19971 = n4886 & n19970;
  assign n19972 = ~n19961 & ~n19971;
  assign n19973 = ~n19949 & n19972;
  assign n19974 = ~n4128 & n19352;
  assign n19975 = ~n4845 & n19974;
  assign n19976 = n5057 & n19975;
  assign n19977 = pi128 & ~n501;
  assign n19978 = n5714 & n19977;
  assign n19979 = n5725 & n19978;
  assign n19980 = ~n1172 & n19979;
  assign n19981 = ~n996 & n19980;
  assign n19982 = ~n2306 & n19981;
  assign n19983 = n3819 & n19982;
  assign n19984 = n3821 & n19983;
  assign n19985 = n5736 & n19984;
  assign n19986 = n19897 & n19985;
  assign n19987 = ~n4003 & n19395;
  assign n19988 = ~n4844 & n19987;
  assign n19989 = ~n4903 & n19988;
  assign n19990 = n4909 & n19989;
  assign n19991 = ~n19986 & ~n19990;
  assign n19992 = ~n19976 & n19991;
  assign n19993 = pi112 & ~n4858;
  assign n19994 = ~n4845 & n19993;
  assign n19995 = ~n4841 & n19994;
  assign n19996 = n4879 & n19995;
  assign n19997 = n4823 & n19996;
  assign n19998 = pi120 & ~n501;
  assign n19999 = n4792 & n19998;
  assign n20000 = n4790 & n19999;
  assign n20001 = n4800 & n20000;
  assign n20002 = ~n996 & n20001;
  assign n20003 = ~n2306 & n20002;
  assign n20004 = n3819 & n20003;
  assign n20005 = n4789 & n20004;
  assign n20006 = n3823 & n20005;
  assign n20007 = n5689 & n20006;
  assign n20008 = n5560 & n20007;
  assign n20009 = n5201 & n20008;
  assign n20010 = ~n5112 & n20009;
  assign n20011 = n5710 & n20010;
  assign n20012 = ~n19997 & ~n20011;
  assign n20013 = n4095 & n19386;
  assign n20014 = n5062 & n20013;
  assign n20015 = n5068 & n20014;
  assign n20016 = n5029 & n20015;
  assign n20017 = ~n5028 & n20016;
  assign n20018 = ~n3940 & n20017;
  assign n20019 = ~n4001 & n20018;
  assign n20020 = ~n4845 & n20019;
  assign n20021 = n5041 & n20020;
  assign n20022 = n5027 & n20021;
  assign n20023 = n1056 & n18169;
  assign n20024 = ~n1208 & n20023;
  assign n20025 = n4920 & n20024;
  assign n20026 = n4925 & n20025;
  assign n20027 = n4932 & n20026;
  assign n20028 = ~n4917 & n20027;
  assign n20029 = ~n1372 & n20028;
  assign n20030 = ~n2243 & n20029;
  assign n20031 = ~n3104 & n20030;
  assign n20032 = ~n3971 & n20031;
  assign n20033 = ~n4003 & n20032;
  assign n20034 = ~n4872 & n20033;
  assign n20035 = ~n4916 & n20034;
  assign n20036 = n4944 & n20035;
  assign n20037 = n4915 & n20036;
  assign n20038 = ~n20022 & ~n20037;
  assign n20039 = n20012 & n20038;
  assign n20040 = n19992 & n20039;
  assign po065 = ~n19973 | ~n20040;
  assign n20042 = n2573 & n18912;
  assign n20043 = n5002 & n20042;
  assign n20044 = n5010 & n20043;
  assign n20045 = n4983 & n20044;
  assign n20046 = ~n4981 & n20045;
  assign n20047 = ~n3066 & n20046;
  assign n20048 = ~n3983 & n20047;
  assign n20049 = ~n4003 & n20048;
  assign n20050 = ~n4024 & n20049;
  assign n20051 = ~n4980 & n20050;
  assign n20052 = n4997 & n20051;
  assign n20053 = n4979 & n20052;
  assign n20054 = pi113 & ~n4858;
  assign n20055 = ~n4845 & n20054;
  assign n20056 = ~n4841 & n20055;
  assign n20057 = n4879 & n20056;
  assign n20058 = n4823 & n20057;
  assign n20059 = pi105 & ~n4648;
  assign n20060 = n5087 & n20059;
  assign n20061 = n5085 & n20060;
  assign n20062 = n5097 & n20061;
  assign n20063 = n4889 & n20062;
  assign n20064 = ~n4887 & n20063;
  assign n20065 = ~n4817 & n20064;
  assign n20066 = ~n4845 & n20065;
  assign n20067 = n4900 & n20066;
  assign n20068 = n4886 & n20067;
  assign n20069 = ~n20058 & ~n20068;
  assign n20070 = ~n20053 & n20069;
  assign n20071 = pi121 & ~n501;
  assign n20072 = n4792 & n20071;
  assign n20073 = n4790 & n20072;
  assign n20074 = n4800 & n20073;
  assign n20075 = ~n996 & n20074;
  assign n20076 = ~n2306 & n20075;
  assign n20077 = n3819 & n20076;
  assign n20078 = n4789 & n20077;
  assign n20079 = n3823 & n20078;
  assign n20080 = n5689 & n20079;
  assign n20081 = n5560 & n20080;
  assign n20082 = n5201 & n20081;
  assign n20083 = ~n5112 & n20082;
  assign n20084 = n5710 & n20083;
  assign n20085 = pi129 & ~n501;
  assign n20086 = n5714 & n20085;
  assign n20087 = n5725 & n20086;
  assign n20088 = ~n1172 & n20087;
  assign n20089 = ~n996 & n20088;
  assign n20090 = ~n2306 & n20089;
  assign n20091 = n3819 & n20090;
  assign n20092 = n3821 & n20091;
  assign n20093 = n5736 & n20092;
  assign n20094 = n19897 & n20093;
  assign n20095 = ~n4003 & n19466;
  assign n20096 = ~n4844 & n20095;
  assign n20097 = ~n4903 & n20096;
  assign n20098 = n4909 & n20097;
  assign n20099 = ~n20094 & ~n20098;
  assign n20100 = ~n20084 & n20099;
  assign n20101 = ~n4128 & n19423;
  assign n20102 = ~n4845 & n20101;
  assign n20103 = n5057 & n20102;
  assign n20104 = n4095 & n19437;
  assign n20105 = n5062 & n20104;
  assign n20106 = n5068 & n20105;
  assign n20107 = n5029 & n20106;
  assign n20108 = ~n5028 & n20107;
  assign n20109 = ~n3940 & n20108;
  assign n20110 = ~n4001 & n20109;
  assign n20111 = ~n4845 & n20110;
  assign n20112 = n5041 & n20111;
  assign n20113 = n5027 & n20112;
  assign n20114 = ~n20103 & ~n20113;
  assign n20115 = n1928 & n18542;
  assign n20116 = n4959 & n20115;
  assign n20117 = n4958 & n20116;
  assign n20118 = ~n4953 & n20117;
  assign n20119 = ~n2242 & n20118;
  assign n20120 = ~n3095 & n20119;
  assign n20121 = ~n3997 & n20120;
  assign n20122 = ~n4003 & n20121;
  assign n20123 = ~n4837 & n20122;
  assign n20124 = ~n4952 & n20123;
  assign n20125 = n4972 & n20124;
  assign n20126 = n4951 & n20125;
  assign n20127 = n1056 & n18181;
  assign n20128 = ~n1208 & n20127;
  assign n20129 = n4920 & n20128;
  assign n20130 = n4925 & n20129;
  assign n20131 = n4932 & n20130;
  assign n20132 = ~n4917 & n20131;
  assign n20133 = ~n1372 & n20132;
  assign n20134 = ~n2243 & n20133;
  assign n20135 = ~n3104 & n20134;
  assign n20136 = ~n3971 & n20135;
  assign n20137 = ~n4003 & n20136;
  assign n20138 = ~n4872 & n20137;
  assign n20139 = ~n4916 & n20138;
  assign n20140 = n4944 & n20139;
  assign n20141 = n4915 & n20140;
  assign n20142 = ~n20126 & ~n20141;
  assign n20143 = n20114 & n20142;
  assign n20144 = n20100 & n20143;
  assign po066 = ~n20070 | ~n20144;
  assign n20146 = n4095 & n19508;
  assign n20147 = n5062 & n20146;
  assign n20148 = n5068 & n20147;
  assign n20149 = n5029 & n20148;
  assign n20150 = ~n5028 & n20149;
  assign n20151 = ~n3940 & n20150;
  assign n20152 = ~n4001 & n20151;
  assign n20153 = ~n4845 & n20152;
  assign n20154 = n5041 & n20153;
  assign n20155 = n5027 & n20154;
  assign n20156 = n1928 & n18580;
  assign n20157 = n4959 & n20156;
  assign n20158 = n4958 & n20157;
  assign n20159 = ~n4953 & n20158;
  assign n20160 = ~n2242 & n20159;
  assign n20161 = ~n3095 & n20160;
  assign n20162 = ~n3997 & n20161;
  assign n20163 = ~n4003 & n20162;
  assign n20164 = ~n4837 & n20163;
  assign n20165 = ~n4952 & n20164;
  assign n20166 = n4972 & n20165;
  assign n20167 = n4951 & n20166;
  assign n20168 = pi122 & ~n501;
  assign n20169 = n4792 & n20168;
  assign n20170 = n4790 & n20169;
  assign n20171 = n4800 & n20170;
  assign n20172 = ~n996 & n20171;
  assign n20173 = ~n2306 & n20172;
  assign n20174 = n3819 & n20173;
  assign n20175 = n4789 & n20174;
  assign n20176 = n3823 & n20175;
  assign n20177 = n5689 & n20176;
  assign n20178 = n5560 & n20177;
  assign n20179 = n5201 & n20178;
  assign n20180 = ~n5112 & n20179;
  assign n20181 = n5710 & n20180;
  assign n20182 = ~n20167 & ~n20181;
  assign n20183 = ~n20155 & n20182;
  assign n20184 = n1056 & n18193;
  assign n20185 = ~n1208 & n20184;
  assign n20186 = n4920 & n20185;
  assign n20187 = n4925 & n20186;
  assign n20188 = n4932 & n20187;
  assign n20189 = ~n4917 & n20188;
  assign n20190 = ~n1372 & n20189;
  assign n20191 = ~n2243 & n20190;
  assign n20192 = ~n3104 & n20191;
  assign n20193 = ~n3971 & n20192;
  assign n20194 = ~n4003 & n20193;
  assign n20195 = ~n4872 & n20194;
  assign n20196 = ~n4916 & n20195;
  assign n20197 = n4944 & n20196;
  assign n20198 = n4915 & n20197;
  assign n20199 = ~n4003 & n19537;
  assign n20200 = ~n4844 & n20199;
  assign n20201 = ~n4903 & n20200;
  assign n20202 = n4909 & n20201;
  assign n20203 = pi130 & ~n501;
  assign n20204 = n5714 & n20203;
  assign n20205 = n5725 & n20204;
  assign n20206 = ~n1172 & n20205;
  assign n20207 = ~n996 & n20206;
  assign n20208 = ~n2306 & n20207;
  assign n20209 = n3819 & n20208;
  assign n20210 = n3821 & n20209;
  assign n20211 = n5736 & n20210;
  assign n20212 = n19897 & n20211;
  assign n20213 = ~n20202 & ~n20212;
  assign n20214 = ~n20198 & n20213;
  assign n20215 = pi114 & ~n4858;
  assign n20216 = ~n4845 & n20215;
  assign n20217 = ~n4841 & n20216;
  assign n20218 = n4879 & n20217;
  assign n20219 = n4823 & n20218;
  assign n20220 = pi106 & ~n4648;
  assign n20221 = n5087 & n20220;
  assign n20222 = n5085 & n20221;
  assign n20223 = n5097 & n20222;
  assign n20224 = n4889 & n20223;
  assign n20225 = ~n4887 & n20224;
  assign n20226 = ~n4817 & n20225;
  assign n20227 = ~n4845 & n20226;
  assign n20228 = n4900 & n20227;
  assign n20229 = n4886 & n20228;
  assign n20230 = ~n20219 & ~n20229;
  assign n20231 = ~n4128 & n19494;
  assign n20232 = ~n4845 & n20231;
  assign n20233 = n5057 & n20232;
  assign n20234 = n2573 & n18971;
  assign n20235 = n5002 & n20234;
  assign n20236 = n5010 & n20235;
  assign n20237 = n4983 & n20236;
  assign n20238 = ~n4981 & n20237;
  assign n20239 = ~n3066 & n20238;
  assign n20240 = ~n3983 & n20239;
  assign n20241 = ~n4003 & n20240;
  assign n20242 = ~n4024 & n20241;
  assign n20243 = ~n4980 & n20242;
  assign n20244 = n4997 & n20243;
  assign n20245 = n4979 & n20244;
  assign n20246 = ~n20233 & ~n20245;
  assign n20247 = n20230 & n20246;
  assign n20248 = n20214 & n20247;
  assign po067 = ~n20183 | ~n20248;
  assign n20250 = n1928 & n18618;
  assign n20251 = n4959 & n20250;
  assign n20252 = n4958 & n20251;
  assign n20253 = ~n4953 & n20252;
  assign n20254 = ~n2242 & n20253;
  assign n20255 = ~n3095 & n20254;
  assign n20256 = ~n3997 & n20255;
  assign n20257 = ~n4003 & n20256;
  assign n20258 = ~n4837 & n20257;
  assign n20259 = ~n4952 & n20258;
  assign n20260 = n4972 & n20259;
  assign n20261 = n4951 & n20260;
  assign n20262 = pi123 & ~n501;
  assign n20263 = n4792 & n20262;
  assign n20264 = n4790 & n20263;
  assign n20265 = n4800 & n20264;
  assign n20266 = ~n996 & n20265;
  assign n20267 = ~n2306 & n20266;
  assign n20268 = n3819 & n20267;
  assign n20269 = n4789 & n20268;
  assign n20270 = n3823 & n20269;
  assign n20271 = n5689 & n20270;
  assign n20272 = n5560 & n20271;
  assign n20273 = n5201 & n20272;
  assign n20274 = ~n5112 & n20273;
  assign n20275 = n5710 & n20274;
  assign n20276 = n4095 & n19579;
  assign n20277 = n5062 & n20276;
  assign n20278 = n5068 & n20277;
  assign n20279 = n5029 & n20278;
  assign n20280 = ~n5028 & n20279;
  assign n20281 = ~n3940 & n20280;
  assign n20282 = ~n4001 & n20281;
  assign n20283 = ~n4845 & n20282;
  assign n20284 = n5041 & n20283;
  assign n20285 = n5027 & n20284;
  assign n20286 = ~n20275 & ~n20285;
  assign n20287 = ~n20261 & n20286;
  assign n20288 = n1056 & n18205;
  assign n20289 = ~n1208 & n20288;
  assign n20290 = n4920 & n20289;
  assign n20291 = n4925 & n20290;
  assign n20292 = n4932 & n20291;
  assign n20293 = ~n4917 & n20292;
  assign n20294 = ~n1372 & n20293;
  assign n20295 = ~n2243 & n20294;
  assign n20296 = ~n3104 & n20295;
  assign n20297 = ~n3971 & n20296;
  assign n20298 = ~n4003 & n20297;
  assign n20299 = ~n4872 & n20298;
  assign n20300 = ~n4916 & n20299;
  assign n20301 = n4944 & n20300;
  assign n20302 = n4915 & n20301;
  assign n20303 = ~n4003 & n19608;
  assign n20304 = ~n4844 & n20303;
  assign n20305 = ~n4903 & n20304;
  assign n20306 = n4909 & n20305;
  assign n20307 = pi131 & ~n501;
  assign n20308 = n5714 & n20307;
  assign n20309 = n5725 & n20308;
  assign n20310 = ~n1172 & n20309;
  assign n20311 = ~n996 & n20310;
  assign n20312 = ~n2306 & n20311;
  assign n20313 = n3819 & n20312;
  assign n20314 = n3821 & n20313;
  assign n20315 = n5736 & n20314;
  assign n20316 = n19897 & n20315;
  assign n20317 = ~n20306 & ~n20316;
  assign n20318 = ~n20302 & n20317;
  assign n20319 = pi115 & ~n4858;
  assign n20320 = ~n4845 & n20319;
  assign n20321 = ~n4841 & n20320;
  assign n20322 = n4879 & n20321;
  assign n20323 = n4823 & n20322;
  assign n20324 = pi107 & ~n4648;
  assign n20325 = n5087 & n20324;
  assign n20326 = n5085 & n20325;
  assign n20327 = n5097 & n20326;
  assign n20328 = n4889 & n20327;
  assign n20329 = ~n4887 & n20328;
  assign n20330 = ~n4817 & n20329;
  assign n20331 = ~n4845 & n20330;
  assign n20332 = n4900 & n20331;
  assign n20333 = n4886 & n20332;
  assign n20334 = ~n20323 & ~n20333;
  assign n20335 = ~n4128 & n19565;
  assign n20336 = ~n4845 & n20335;
  assign n20337 = n5057 & n20336;
  assign n20338 = n2573 & n19030;
  assign n20339 = n5002 & n20338;
  assign n20340 = n5010 & n20339;
  assign n20341 = n4983 & n20340;
  assign n20342 = ~n4981 & n20341;
  assign n20343 = ~n3066 & n20342;
  assign n20344 = ~n3983 & n20343;
  assign n20345 = ~n4003 & n20344;
  assign n20346 = ~n4024 & n20345;
  assign n20347 = ~n4980 & n20346;
  assign n20348 = n4997 & n20347;
  assign n20349 = n4979 & n20348;
  assign n20350 = ~n20337 & ~n20349;
  assign n20351 = n20334 & n20350;
  assign n20352 = n20318 & n20351;
  assign po068 = ~n20287 | ~n20352;
  assign n20354 = n1928 & n18656;
  assign n20355 = n4959 & n20354;
  assign n20356 = n4958 & n20355;
  assign n20357 = ~n4953 & n20356;
  assign n20358 = ~n2242 & n20357;
  assign n20359 = ~n3095 & n20358;
  assign n20360 = ~n3997 & n20359;
  assign n20361 = ~n4003 & n20360;
  assign n20362 = ~n4837 & n20361;
  assign n20363 = ~n4952 & n20362;
  assign n20364 = n4972 & n20363;
  assign n20365 = n4951 & n20364;
  assign n20366 = pi124 & ~n501;
  assign n20367 = n4792 & n20366;
  assign n20368 = n4790 & n20367;
  assign n20369 = n4800 & n20368;
  assign n20370 = ~n996 & n20369;
  assign n20371 = ~n2306 & n20370;
  assign n20372 = n3819 & n20371;
  assign n20373 = n4789 & n20372;
  assign n20374 = n3823 & n20373;
  assign n20375 = n5689 & n20374;
  assign n20376 = n5560 & n20375;
  assign n20377 = n5201 & n20376;
  assign n20378 = ~n5112 & n20377;
  assign n20379 = n5710 & n20378;
  assign n20380 = n4095 & n19650;
  assign n20381 = n5062 & n20380;
  assign n20382 = n5068 & n20381;
  assign n20383 = n5029 & n20382;
  assign n20384 = ~n5028 & n20383;
  assign n20385 = ~n3940 & n20384;
  assign n20386 = ~n4001 & n20385;
  assign n20387 = ~n4845 & n20386;
  assign n20388 = n5041 & n20387;
  assign n20389 = n5027 & n20388;
  assign n20390 = ~n20379 & ~n20389;
  assign n20391 = ~n20365 & n20390;
  assign n20392 = n1056 & n18217;
  assign n20393 = ~n1208 & n20392;
  assign n20394 = n4920 & n20393;
  assign n20395 = n4925 & n20394;
  assign n20396 = n4932 & n20395;
  assign n20397 = ~n4917 & n20396;
  assign n20398 = ~n1372 & n20397;
  assign n20399 = ~n2243 & n20398;
  assign n20400 = ~n3104 & n20399;
  assign n20401 = ~n3971 & n20400;
  assign n20402 = ~n4003 & n20401;
  assign n20403 = ~n4872 & n20402;
  assign n20404 = ~n4916 & n20403;
  assign n20405 = n4944 & n20404;
  assign n20406 = n4915 & n20405;
  assign n20407 = ~n4003 & n19679;
  assign n20408 = ~n4844 & n20407;
  assign n20409 = ~n4903 & n20408;
  assign n20410 = n4909 & n20409;
  assign n20411 = pi132 & ~n501;
  assign n20412 = n5714 & n20411;
  assign n20413 = n5725 & n20412;
  assign n20414 = ~n1172 & n20413;
  assign n20415 = ~n996 & n20414;
  assign n20416 = ~n2306 & n20415;
  assign n20417 = n3819 & n20416;
  assign n20418 = n3821 & n20417;
  assign n20419 = n5736 & n20418;
  assign n20420 = n19897 & n20419;
  assign n20421 = ~n20410 & ~n20420;
  assign n20422 = ~n20406 & n20421;
  assign n20423 = pi116 & ~n4858;
  assign n20424 = ~n4845 & n20423;
  assign n20425 = ~n4841 & n20424;
  assign n20426 = n4879 & n20425;
  assign n20427 = n4823 & n20426;
  assign n20428 = pi108 & ~n4648;
  assign n20429 = n5087 & n20428;
  assign n20430 = n5085 & n20429;
  assign n20431 = n5097 & n20430;
  assign n20432 = n4889 & n20431;
  assign n20433 = ~n4887 & n20432;
  assign n20434 = ~n4817 & n20433;
  assign n20435 = ~n4845 & n20434;
  assign n20436 = n4900 & n20435;
  assign n20437 = n4886 & n20436;
  assign n20438 = ~n20427 & ~n20437;
  assign n20439 = ~n4128 & n19636;
  assign n20440 = ~n4845 & n20439;
  assign n20441 = n5057 & n20440;
  assign n20442 = n2573 & n19089;
  assign n20443 = n5002 & n20442;
  assign n20444 = n5010 & n20443;
  assign n20445 = n4983 & n20444;
  assign n20446 = ~n4981 & n20445;
  assign n20447 = ~n3066 & n20446;
  assign n20448 = ~n3983 & n20447;
  assign n20449 = ~n4003 & n20448;
  assign n20450 = ~n4024 & n20449;
  assign n20451 = ~n4980 & n20450;
  assign n20452 = n4997 & n20451;
  assign n20453 = n4979 & n20452;
  assign n20454 = ~n20441 & ~n20453;
  assign n20455 = n20438 & n20454;
  assign n20456 = n20422 & n20455;
  assign po069 = ~n20391 | ~n20456;
  assign n20458 = n1928 & n18694;
  assign n20459 = n4959 & n20458;
  assign n20460 = n4958 & n20459;
  assign n20461 = ~n4953 & n20460;
  assign n20462 = ~n2242 & n20461;
  assign n20463 = ~n3095 & n20462;
  assign n20464 = ~n3997 & n20463;
  assign n20465 = ~n4003 & n20464;
  assign n20466 = ~n4837 & n20465;
  assign n20467 = ~n4952 & n20466;
  assign n20468 = n4972 & n20467;
  assign n20469 = n4951 & n20468;
  assign n20470 = pi125 & ~n501;
  assign n20471 = n4792 & n20470;
  assign n20472 = n4790 & n20471;
  assign n20473 = n4800 & n20472;
  assign n20474 = ~n996 & n20473;
  assign n20475 = ~n2306 & n20474;
  assign n20476 = n3819 & n20475;
  assign n20477 = n4789 & n20476;
  assign n20478 = n3823 & n20477;
  assign n20479 = n5689 & n20478;
  assign n20480 = n5560 & n20479;
  assign n20481 = n5201 & n20480;
  assign n20482 = ~n5112 & n20481;
  assign n20483 = n5710 & n20482;
  assign n20484 = n4095 & n19721;
  assign n20485 = n5062 & n20484;
  assign n20486 = n5068 & n20485;
  assign n20487 = n5029 & n20486;
  assign n20488 = ~n5028 & n20487;
  assign n20489 = ~n3940 & n20488;
  assign n20490 = ~n4001 & n20489;
  assign n20491 = ~n4845 & n20490;
  assign n20492 = n5041 & n20491;
  assign n20493 = n5027 & n20492;
  assign n20494 = ~n20483 & ~n20493;
  assign n20495 = ~n20469 & n20494;
  assign n20496 = n1056 & n18229;
  assign n20497 = ~n1208 & n20496;
  assign n20498 = n4920 & n20497;
  assign n20499 = n4925 & n20498;
  assign n20500 = n4932 & n20499;
  assign n20501 = ~n4917 & n20500;
  assign n20502 = ~n1372 & n20501;
  assign n20503 = ~n2243 & n20502;
  assign n20504 = ~n3104 & n20503;
  assign n20505 = ~n3971 & n20504;
  assign n20506 = ~n4003 & n20505;
  assign n20507 = ~n4872 & n20506;
  assign n20508 = ~n4916 & n20507;
  assign n20509 = n4944 & n20508;
  assign n20510 = n4915 & n20509;
  assign n20511 = ~n4003 & n19750;
  assign n20512 = ~n4844 & n20511;
  assign n20513 = ~n4903 & n20512;
  assign n20514 = n4909 & n20513;
  assign n20515 = pi133 & ~n501;
  assign n20516 = n5714 & n20515;
  assign n20517 = n5725 & n20516;
  assign n20518 = ~n1172 & n20517;
  assign n20519 = ~n996 & n20518;
  assign n20520 = ~n2306 & n20519;
  assign n20521 = n3819 & n20520;
  assign n20522 = n3821 & n20521;
  assign n20523 = n5736 & n20522;
  assign n20524 = n19897 & n20523;
  assign n20525 = ~n20514 & ~n20524;
  assign n20526 = ~n20510 & n20525;
  assign n20527 = pi117 & ~n4858;
  assign n20528 = ~n4845 & n20527;
  assign n20529 = ~n4841 & n20528;
  assign n20530 = n4879 & n20529;
  assign n20531 = n4823 & n20530;
  assign n20532 = pi109 & ~n4648;
  assign n20533 = n5087 & n20532;
  assign n20534 = n5085 & n20533;
  assign n20535 = n5097 & n20534;
  assign n20536 = n4889 & n20535;
  assign n20537 = ~n4887 & n20536;
  assign n20538 = ~n4817 & n20537;
  assign n20539 = ~n4845 & n20538;
  assign n20540 = n4900 & n20539;
  assign n20541 = n4886 & n20540;
  assign n20542 = ~n20531 & ~n20541;
  assign n20543 = ~n4128 & n19707;
  assign n20544 = ~n4845 & n20543;
  assign n20545 = n5057 & n20544;
  assign n20546 = n2573 & n19148;
  assign n20547 = n5002 & n20546;
  assign n20548 = n5010 & n20547;
  assign n20549 = n4983 & n20548;
  assign n20550 = ~n4981 & n20549;
  assign n20551 = ~n3066 & n20550;
  assign n20552 = ~n3983 & n20551;
  assign n20553 = ~n4003 & n20552;
  assign n20554 = ~n4024 & n20553;
  assign n20555 = ~n4980 & n20554;
  assign n20556 = n4997 & n20555;
  assign n20557 = n4979 & n20556;
  assign n20558 = ~n20545 & ~n20557;
  assign n20559 = n20542 & n20558;
  assign n20560 = n20526 & n20559;
  assign po070 = ~n20495 | ~n20560;
  assign n20562 = n1928 & n18732;
  assign n20563 = n4959 & n20562;
  assign n20564 = n4958 & n20563;
  assign n20565 = ~n4953 & n20564;
  assign n20566 = ~n2242 & n20565;
  assign n20567 = ~n3095 & n20566;
  assign n20568 = ~n3997 & n20567;
  assign n20569 = ~n4003 & n20568;
  assign n20570 = ~n4837 & n20569;
  assign n20571 = ~n4952 & n20570;
  assign n20572 = n4972 & n20571;
  assign n20573 = n4951 & n20572;
  assign n20574 = pi126 & ~n501;
  assign n20575 = n4792 & n20574;
  assign n20576 = n4790 & n20575;
  assign n20577 = n4800 & n20576;
  assign n20578 = ~n996 & n20577;
  assign n20579 = ~n2306 & n20578;
  assign n20580 = n3819 & n20579;
  assign n20581 = n4789 & n20580;
  assign n20582 = n3823 & n20581;
  assign n20583 = n5689 & n20582;
  assign n20584 = n5560 & n20583;
  assign n20585 = n5201 & n20584;
  assign n20586 = ~n5112 & n20585;
  assign n20587 = n5710 & n20586;
  assign n20588 = n4095 & n19792;
  assign n20589 = n5062 & n20588;
  assign n20590 = n5068 & n20589;
  assign n20591 = n5029 & n20590;
  assign n20592 = ~n5028 & n20591;
  assign n20593 = ~n3940 & n20592;
  assign n20594 = ~n4001 & n20593;
  assign n20595 = ~n4845 & n20594;
  assign n20596 = n5041 & n20595;
  assign n20597 = n5027 & n20596;
  assign n20598 = ~n20587 & ~n20597;
  assign n20599 = ~n20573 & n20598;
  assign n20600 = n1056 & n18241;
  assign n20601 = ~n1208 & n20600;
  assign n20602 = n4920 & n20601;
  assign n20603 = n4925 & n20602;
  assign n20604 = n4932 & n20603;
  assign n20605 = ~n4917 & n20604;
  assign n20606 = ~n1372 & n20605;
  assign n20607 = ~n2243 & n20606;
  assign n20608 = ~n3104 & n20607;
  assign n20609 = ~n3971 & n20608;
  assign n20610 = ~n4003 & n20609;
  assign n20611 = ~n4872 & n20610;
  assign n20612 = ~n4916 & n20611;
  assign n20613 = n4944 & n20612;
  assign n20614 = n4915 & n20613;
  assign n20615 = ~n4003 & n19821;
  assign n20616 = ~n4844 & n20615;
  assign n20617 = ~n4903 & n20616;
  assign n20618 = n4909 & n20617;
  assign n20619 = pi134 & ~n501;
  assign n20620 = n5714 & n20619;
  assign n20621 = n5725 & n20620;
  assign n20622 = ~n1172 & n20621;
  assign n20623 = ~n996 & n20622;
  assign n20624 = ~n2306 & n20623;
  assign n20625 = n3819 & n20624;
  assign n20626 = n3821 & n20625;
  assign n20627 = n5736 & n20626;
  assign n20628 = n19897 & n20627;
  assign n20629 = ~n20618 & ~n20628;
  assign n20630 = ~n20614 & n20629;
  assign n20631 = pi118 & ~n4858;
  assign n20632 = ~n4845 & n20631;
  assign n20633 = ~n4841 & n20632;
  assign n20634 = n4879 & n20633;
  assign n20635 = n4823 & n20634;
  assign n20636 = pi110 & ~n4648;
  assign n20637 = n5087 & n20636;
  assign n20638 = n5085 & n20637;
  assign n20639 = n5097 & n20638;
  assign n20640 = n4889 & n20639;
  assign n20641 = ~n4887 & n20640;
  assign n20642 = ~n4817 & n20641;
  assign n20643 = ~n4845 & n20642;
  assign n20644 = n4900 & n20643;
  assign n20645 = n4886 & n20644;
  assign n20646 = ~n20635 & ~n20645;
  assign n20647 = ~n4128 & n19778;
  assign n20648 = ~n4845 & n20647;
  assign n20649 = n5057 & n20648;
  assign n20650 = n2573 & n19207;
  assign n20651 = n5002 & n20650;
  assign n20652 = n5010 & n20651;
  assign n20653 = n4983 & n20652;
  assign n20654 = ~n4981 & n20653;
  assign n20655 = ~n3066 & n20654;
  assign n20656 = ~n3983 & n20655;
  assign n20657 = ~n4003 & n20656;
  assign n20658 = ~n4024 & n20657;
  assign n20659 = ~n4980 & n20658;
  assign n20660 = n4997 & n20659;
  assign n20661 = n4979 & n20660;
  assign n20662 = ~n20649 & ~n20661;
  assign n20663 = n20646 & n20662;
  assign n20664 = n20630 & n20663;
  assign po071 = ~n20599 | ~n20664;
  assign n20666 = n5837 & n18466;
  assign n20667 = n5839 & n20666;
  assign n20668 = n5836 & n20667;
  assign n20669 = ~n5834 & n20668;
  assign n20670 = ~n2242 & n20669;
  assign n20671 = ~n3095 & n20670;
  assign n20672 = ~n3997 & n20671;
  assign n20673 = ~n4003 & n20672;
  assign n20674 = ~n4837 & n20673;
  assign n20675 = ~n5822 & n20674;
  assign n20676 = ~n5833 & n20675;
  assign n20677 = n5856 & n20676;
  assign n20678 = n5832 & n20677;
  assign n20679 = pi087 & ~n3340;
  assign n20680 = ~n3341 & n20679;
  assign n20681 = ~n3339 & n20680;
  assign n20682 = ~n3524 & n20681;
  assign n20683 = n4097 & n20682;
  assign n20684 = ~n3373 & ~n3679;
  assign n20685 = n3433 & n20684;
  assign n20686 = n4104 & n20685;
  assign n20687 = n20683 & n20686;
  assign n20688 = n5925 & n20687;
  assign n20689 = ~n5924 & n20688;
  assign n20690 = ~n3940 & n20689;
  assign n20691 = ~n4001 & n20690;
  assign n20692 = ~n5043 & n20691;
  assign n20693 = ~n5923 & n20692;
  assign n20694 = n5941 & n20693;
  assign n20695 = n5922 & n20694;
  assign n20696 = pi103 & ~n4677;
  assign n20697 = n4737 & n20696;
  assign n20698 = n4491 & n20697;
  assign n20699 = n4891 & n20698;
  assign n20700 = n5986 & n20699;
  assign n20701 = ~n5985 & n20700;
  assign n20702 = ~n4817 & n20701;
  assign n20703 = ~n4902 & n20702;
  assign n20704 = ~n5923 & n20703;
  assign n20705 = n5999 & n20704;
  assign n20706 = n5984 & n20705;
  assign n20707 = ~n20695 & ~n20706;
  assign n20708 = ~n20678 & n20707;
  assign n20709 = pi143 & ~n501;
  assign n20710 = n5713 & n20709;
  assign n20711 = n6138 & n20710;
  assign n20712 = n6147 & n20711;
  assign n20713 = ~n1172 & n20712;
  assign n20714 = ~n996 & n20713;
  assign n20715 = ~n2306 & n20714;
  assign n20716 = n3819 & n20715;
  assign n20717 = n3821 & n20716;
  assign n20718 = n6183 & n20717;
  assign n20719 = n19897 & n20718;
  assign n20720 = ~n6137 & n20719;
  assign n20721 = n6193 & n20720;
  assign n20722 = n6134 & n20721;
  assign n20723 = ~n5911 & n19884;
  assign n20724 = ~n5909 & n20723;
  assign n20725 = n5916 & n20724;
  assign n20726 = pi135 & ~n501;
  assign n20727 = n6687 & n20726;
  assign n20728 = n6685 & n20727;
  assign n20729 = n6692 & n20728;
  assign n20730 = n6683 & n20729;
  assign n20731 = ~n1172 & n20730;
  assign n20732 = ~n1054 & n20731;
  assign n20733 = ~n996 & n20732;
  assign n20734 = n6698 & n20733;
  assign n20735 = n6677 & n20734;
  assign n20736 = n6707 & n20735;
  assign n20737 = n6711 & n20736;
  assign n20738 = n6676 & n20737;
  assign n20739 = n6284 & n20738;
  assign n20740 = ~n20725 & ~n20739;
  assign n20741 = ~n20722 & n20740;
  assign n20742 = ~n5058 & n19931;
  assign n20743 = ~n5923 & n20742;
  assign n20744 = n5966 & n20743;
  assign n20745 = ~n4881 & n19926;
  assign n20746 = ~n5923 & n20745;
  assign n20747 = n6025 & n20746;
  assign n20748 = n6021 & n20747;
  assign n20749 = ~n20744 & ~n20748;
  assign n20750 = n20741 & n20749;
  assign n20751 = pi039 & ~n1144;
  assign n20752 = ~n1115 & n20751;
  assign n20753 = n1056 & n20752;
  assign n20754 = ~n1208 & n20753;
  assign n20755 = n4920 & n20754;
  assign n20756 = n5873 & n20755;
  assign n20757 = n4932 & n20756;
  assign n20758 = ~n5865 & n20757;
  assign n20759 = ~n1372 & n20758;
  assign n20760 = ~n2243 & n20759;
  assign n20761 = ~n3104 & n20760;
  assign n20762 = ~n3971 & n20761;
  assign n20763 = ~n4003 & n20762;
  assign n20764 = ~n4872 & n20763;
  assign n20765 = ~n5801 & n20764;
  assign n20766 = ~n5864 & n20765;
  assign n20767 = n5891 & n20766;
  assign n20768 = n5863 & n20767;
  assign n20769 = ~n5141 & n6036;
  assign n20770 = pi119 & ~n5523;
  assign n20771 = ~n5172 & ~n5524;
  assign n20772 = n20770 & n20771;
  assign n20773 = ~n5522 & n20772;
  assign n20774 = ~n5598 & n20773;
  assign n20775 = n6068 & n20774;
  assign n20776 = n6066 & n20775;
  assign n20777 = ~n5197 & ~n5318;
  assign n20778 = ~n5498 & n20777;
  assign n20779 = n6075 & n20778;
  assign n20780 = n20776 & n20779;
  assign n20781 = n20769 & n20780;
  assign n20782 = ~n6035 & n20781;
  assign n20783 = ~n5808 & n20782;
  assign n20784 = ~n5923 & n20783;
  assign n20785 = n6054 & n20784;
  assign n20786 = n6034 & n20785;
  assign n20787 = ~n20768 & ~n20786;
  assign n20788 = pi071 & ~n2659;
  assign n20789 = ~n2660 & n20788;
  assign n20790 = ~n2658 & n20789;
  assign n20791 = ~n2363 & n20790;
  assign n20792 = n2633 & n20791;
  assign n20793 = n3977 & n20792;
  assign n20794 = n5771 & n20793;
  assign n20795 = ~n5770 & n20794;
  assign n20796 = ~n3066 & n20795;
  assign n20797 = ~n3983 & n20796;
  assign n20798 = ~n4003 & n20797;
  assign n20799 = ~n4024 & n20798;
  assign n20800 = ~n4999 & n20799;
  assign n20801 = ~n5751 & n20800;
  assign n20802 = n5825 & n20801;
  assign n20803 = n5750 & n20802;
  assign n20804 = pi127 & ~n5769;
  assign n20805 = ~n5923 & n20804;
  assign n20806 = ~n5958 & n20805;
  assign n20807 = n6112 & n20806;
  assign n20808 = n6095 & n20807;
  assign n20809 = ~n20803 & ~n20808;
  assign n20810 = n20787 & n20809;
  assign n20811 = n20750 & n20810;
  assign po072 = ~n20708 | ~n20811;
  assign n20813 = pi040 & ~n1144;
  assign n20814 = ~n1115 & n20813;
  assign n20815 = n1056 & n20814;
  assign n20816 = ~n1208 & n20815;
  assign n20817 = n4920 & n20816;
  assign n20818 = n5873 & n20817;
  assign n20819 = n4932 & n20818;
  assign n20820 = ~n5865 & n20819;
  assign n20821 = ~n1372 & n20820;
  assign n20822 = ~n2243 & n20821;
  assign n20823 = ~n3104 & n20822;
  assign n20824 = ~n3971 & n20823;
  assign n20825 = ~n4003 & n20824;
  assign n20826 = ~n4872 & n20825;
  assign n20827 = ~n5801 & n20826;
  assign n20828 = ~n5864 & n20827;
  assign n20829 = n5891 & n20828;
  assign n20830 = n5863 & n20829;
  assign n20831 = n5837 & n18504;
  assign n20832 = n5839 & n20831;
  assign n20833 = n5836 & n20832;
  assign n20834 = ~n5834 & n20833;
  assign n20835 = ~n2242 & n20834;
  assign n20836 = ~n3095 & n20835;
  assign n20837 = ~n3997 & n20836;
  assign n20838 = ~n4003 & n20837;
  assign n20839 = ~n4837 & n20838;
  assign n20840 = ~n5822 & n20839;
  assign n20841 = ~n5833 & n20840;
  assign n20842 = n5856 & n20841;
  assign n20843 = n5832 & n20842;
  assign n20844 = pi104 & ~n4677;
  assign n20845 = n4737 & n20844;
  assign n20846 = n4491 & n20845;
  assign n20847 = n4891 & n20846;
  assign n20848 = n5986 & n20847;
  assign n20849 = ~n5985 & n20848;
  assign n20850 = ~n4817 & n20849;
  assign n20851 = ~n4902 & n20850;
  assign n20852 = ~n5923 & n20851;
  assign n20853 = n5999 & n20852;
  assign n20854 = n5984 & n20853;
  assign n20855 = ~n20843 & ~n20854;
  assign n20856 = ~n20830 & n20855;
  assign n20857 = ~n5058 & n19974;
  assign n20858 = ~n5923 & n20857;
  assign n20859 = n5966 & n20858;
  assign n20860 = ~n5911 & n19988;
  assign n20861 = ~n5909 & n20860;
  assign n20862 = n5916 & n20861;
  assign n20863 = pi136 & ~n501;
  assign n20864 = n6687 & n20863;
  assign n20865 = n6685 & n20864;
  assign n20866 = n6692 & n20865;
  assign n20867 = n6683 & n20866;
  assign n20868 = ~n1172 & n20867;
  assign n20869 = ~n1054 & n20868;
  assign n20870 = ~n996 & n20869;
  assign n20871 = n6698 & n20870;
  assign n20872 = n6677 & n20871;
  assign n20873 = n6707 & n20872;
  assign n20874 = n6711 & n20873;
  assign n20875 = n6676 & n20874;
  assign n20876 = n6284 & n20875;
  assign n20877 = ~n20862 & ~n20876;
  assign n20878 = ~n20859 & n20877;
  assign n20879 = ~n4881 & n19993;
  assign n20880 = ~n5923 & n20879;
  assign n20881 = n6025 & n20880;
  assign n20882 = n6021 & n20881;
  assign n20883 = pi144 & ~n501;
  assign n20884 = n5713 & n20883;
  assign n20885 = n6138 & n20884;
  assign n20886 = n6147 & n20885;
  assign n20887 = ~n1172 & n20886;
  assign n20888 = ~n996 & n20887;
  assign n20889 = ~n2306 & n20888;
  assign n20890 = n3819 & n20889;
  assign n20891 = n3821 & n20890;
  assign n20892 = n6183 & n20891;
  assign n20893 = n19897 & n20892;
  assign n20894 = ~n6137 & n20893;
  assign n20895 = n6193 & n20894;
  assign n20896 = n6134 & n20895;
  assign n20897 = ~n20882 & ~n20896;
  assign n20898 = n20878 & n20897;
  assign n20899 = pi120 & ~n5598;
  assign n20900 = n6068 & n20899;
  assign n20901 = n6066 & n20900;
  assign n20902 = n6076 & n20901;
  assign n20903 = n6038 & n20902;
  assign n20904 = ~n6035 & n20903;
  assign n20905 = ~n5808 & n20904;
  assign n20906 = ~n5923 & n20905;
  assign n20907 = n6054 & n20906;
  assign n20908 = n6034 & n20907;
  assign n20909 = n5948 & n20014;
  assign n20910 = n5925 & n20909;
  assign n20911 = ~n5924 & n20910;
  assign n20912 = ~n3940 & n20911;
  assign n20913 = ~n4001 & n20912;
  assign n20914 = ~n5043 & n20913;
  assign n20915 = ~n5923 & n20914;
  assign n20916 = n5941 & n20915;
  assign n20917 = n5922 & n20916;
  assign n20918 = ~n20908 & ~n20917;
  assign n20919 = pi128 & ~n5769;
  assign n20920 = ~n5923 & n20919;
  assign n20921 = ~n5958 & n20920;
  assign n20922 = n6112 & n20921;
  assign n20923 = n6095 & n20922;
  assign n20924 = n5897 & n19939;
  assign n20925 = n5771 & n20924;
  assign n20926 = ~n5770 & n20925;
  assign n20927 = ~n3066 & n20926;
  assign n20928 = ~n3983 & n20927;
  assign n20929 = ~n4003 & n20928;
  assign n20930 = ~n4024 & n20929;
  assign n20931 = ~n4999 & n20930;
  assign n20932 = ~n5751 & n20931;
  assign n20933 = n5825 & n20932;
  assign n20934 = n5750 & n20933;
  assign n20935 = ~n20923 & ~n20934;
  assign n20936 = n20918 & n20935;
  assign n20937 = n20898 & n20936;
  assign po073 = ~n20856 | ~n20937;
  assign n20939 = n5897 & n20043;
  assign n20940 = n5771 & n20939;
  assign n20941 = ~n5770 & n20940;
  assign n20942 = ~n3066 & n20941;
  assign n20943 = ~n3983 & n20942;
  assign n20944 = ~n4003 & n20943;
  assign n20945 = ~n4024 & n20944;
  assign n20946 = ~n4999 & n20945;
  assign n20947 = ~n5751 & n20946;
  assign n20948 = n5825 & n20947;
  assign n20949 = n5750 & n20948;
  assign n20950 = n5837 & n18542;
  assign n20951 = n5839 & n20950;
  assign n20952 = n5836 & n20951;
  assign n20953 = ~n5834 & n20952;
  assign n20954 = ~n2242 & n20953;
  assign n20955 = ~n3095 & n20954;
  assign n20956 = ~n3997 & n20955;
  assign n20957 = ~n4003 & n20956;
  assign n20958 = ~n4837 & n20957;
  assign n20959 = ~n5822 & n20958;
  assign n20960 = ~n5833 & n20959;
  assign n20961 = n5856 & n20960;
  assign n20962 = n5832 & n20961;
  assign n20963 = pi041 & ~n1144;
  assign n20964 = ~n1115 & n20963;
  assign n20965 = n1056 & n20964;
  assign n20966 = ~n1208 & n20965;
  assign n20967 = n4920 & n20966;
  assign n20968 = n5873 & n20967;
  assign n20969 = n4932 & n20968;
  assign n20970 = ~n5865 & n20969;
  assign n20971 = ~n1372 & n20970;
  assign n20972 = ~n2243 & n20971;
  assign n20973 = ~n3104 & n20972;
  assign n20974 = ~n3971 & n20973;
  assign n20975 = ~n4003 & n20974;
  assign n20976 = ~n4872 & n20975;
  assign n20977 = ~n5801 & n20976;
  assign n20978 = ~n5864 & n20977;
  assign n20979 = n5891 & n20978;
  assign n20980 = n5863 & n20979;
  assign n20981 = ~n20962 & ~n20980;
  assign n20982 = ~n20949 & n20981;
  assign n20983 = ~n5058 & n20101;
  assign n20984 = ~n5923 & n20983;
  assign n20985 = n5966 & n20984;
  assign n20986 = ~n5911 & n20096;
  assign n20987 = ~n5909 & n20986;
  assign n20988 = n5916 & n20987;
  assign n20989 = pi137 & ~n501;
  assign n20990 = n6687 & n20989;
  assign n20991 = n6685 & n20990;
  assign n20992 = n6692 & n20991;
  assign n20993 = n6683 & n20992;
  assign n20994 = ~n1172 & n20993;
  assign n20995 = ~n1054 & n20994;
  assign n20996 = ~n996 & n20995;
  assign n20997 = n6698 & n20996;
  assign n20998 = n6677 & n20997;
  assign n20999 = n6707 & n20998;
  assign n21000 = n6711 & n20999;
  assign n21001 = n6676 & n21000;
  assign n21002 = n6284 & n21001;
  assign n21003 = ~n20988 & ~n21002;
  assign n21004 = ~n20985 & n21003;
  assign n21005 = ~n4881 & n20054;
  assign n21006 = ~n5923 & n21005;
  assign n21007 = n6025 & n21006;
  assign n21008 = n6021 & n21007;
  assign n21009 = pi145 & ~n501;
  assign n21010 = n5713 & n21009;
  assign n21011 = n6138 & n21010;
  assign n21012 = n6147 & n21011;
  assign n21013 = ~n1172 & n21012;
  assign n21014 = ~n996 & n21013;
  assign n21015 = ~n2306 & n21014;
  assign n21016 = n3819 & n21015;
  assign n21017 = n3821 & n21016;
  assign n21018 = n6183 & n21017;
  assign n21019 = n19897 & n21018;
  assign n21020 = ~n6137 & n21019;
  assign n21021 = n6193 & n21020;
  assign n21022 = n6134 & n21021;
  assign n21023 = ~n21008 & ~n21022;
  assign n21024 = n21004 & n21023;
  assign n21025 = pi121 & ~n5598;
  assign n21026 = n6068 & n21025;
  assign n21027 = n6066 & n21026;
  assign n21028 = n6076 & n21027;
  assign n21029 = n6038 & n21028;
  assign n21030 = ~n6035 & n21029;
  assign n21031 = ~n5808 & n21030;
  assign n21032 = ~n5923 & n21031;
  assign n21033 = n6054 & n21032;
  assign n21034 = n6034 & n21033;
  assign n21035 = pi105 & ~n4677;
  assign n21036 = n4737 & n21035;
  assign n21037 = n4491 & n21036;
  assign n21038 = n4891 & n21037;
  assign n21039 = n5986 & n21038;
  assign n21040 = ~n5985 & n21039;
  assign n21041 = ~n4817 & n21040;
  assign n21042 = ~n4902 & n21041;
  assign n21043 = ~n5923 & n21042;
  assign n21044 = n5999 & n21043;
  assign n21045 = n5984 & n21044;
  assign n21046 = ~n21034 & ~n21045;
  assign n21047 = n5948 & n20105;
  assign n21048 = n5925 & n21047;
  assign n21049 = ~n5924 & n21048;
  assign n21050 = ~n3940 & n21049;
  assign n21051 = ~n4001 & n21050;
  assign n21052 = ~n5043 & n21051;
  assign n21053 = ~n5923 & n21052;
  assign n21054 = n5941 & n21053;
  assign n21055 = n5922 & n21054;
  assign n21056 = pi129 & ~n5769;
  assign n21057 = ~n5923 & n21056;
  assign n21058 = ~n5958 & n21057;
  assign n21059 = n6112 & n21058;
  assign n21060 = n6095 & n21059;
  assign n21061 = ~n21055 & ~n21060;
  assign n21062 = n21046 & n21061;
  assign n21063 = n21024 & n21062;
  assign po074 = ~n20982 | ~n21063;
  assign n21065 = n5897 & n20235;
  assign n21066 = n5771 & n21065;
  assign n21067 = ~n5770 & n21066;
  assign n21068 = ~n3066 & n21067;
  assign n21069 = ~n3983 & n21068;
  assign n21070 = ~n4003 & n21069;
  assign n21071 = ~n4024 & n21070;
  assign n21072 = ~n4999 & n21071;
  assign n21073 = ~n5751 & n21072;
  assign n21074 = n5825 & n21073;
  assign n21075 = n5750 & n21074;
  assign n21076 = n5837 & n18580;
  assign n21077 = n5839 & n21076;
  assign n21078 = n5836 & n21077;
  assign n21079 = ~n5834 & n21078;
  assign n21080 = ~n2242 & n21079;
  assign n21081 = ~n3095 & n21080;
  assign n21082 = ~n3997 & n21081;
  assign n21083 = ~n4003 & n21082;
  assign n21084 = ~n4837 & n21083;
  assign n21085 = ~n5822 & n21084;
  assign n21086 = ~n5833 & n21085;
  assign n21087 = n5856 & n21086;
  assign n21088 = n5832 & n21087;
  assign n21089 = pi042 & ~n1144;
  assign n21090 = ~n1115 & n21089;
  assign n21091 = n1056 & n21090;
  assign n21092 = ~n1208 & n21091;
  assign n21093 = n4920 & n21092;
  assign n21094 = n5873 & n21093;
  assign n21095 = n4932 & n21094;
  assign n21096 = ~n5865 & n21095;
  assign n21097 = ~n1372 & n21096;
  assign n21098 = ~n2243 & n21097;
  assign n21099 = ~n3104 & n21098;
  assign n21100 = ~n3971 & n21099;
  assign n21101 = ~n4003 & n21100;
  assign n21102 = ~n4872 & n21101;
  assign n21103 = ~n5801 & n21102;
  assign n21104 = ~n5864 & n21103;
  assign n21105 = n5891 & n21104;
  assign n21106 = n5863 & n21105;
  assign n21107 = ~n21088 & ~n21106;
  assign n21108 = ~n21075 & n21107;
  assign n21109 = ~n5058 & n20231;
  assign n21110 = ~n5923 & n21109;
  assign n21111 = n5966 & n21110;
  assign n21112 = ~n5911 & n20200;
  assign n21113 = ~n5909 & n21112;
  assign n21114 = n5916 & n21113;
  assign n21115 = pi138 & ~n501;
  assign n21116 = n6687 & n21115;
  assign n21117 = n6685 & n21116;
  assign n21118 = n6692 & n21117;
  assign n21119 = n6683 & n21118;
  assign n21120 = ~n1172 & n21119;
  assign n21121 = ~n1054 & n21120;
  assign n21122 = ~n996 & n21121;
  assign n21123 = n6698 & n21122;
  assign n21124 = n6677 & n21123;
  assign n21125 = n6707 & n21124;
  assign n21126 = n6711 & n21125;
  assign n21127 = n6676 & n21126;
  assign n21128 = n6284 & n21127;
  assign n21129 = ~n21114 & ~n21128;
  assign n21130 = ~n21111 & n21129;
  assign n21131 = ~n4881 & n20215;
  assign n21132 = ~n5923 & n21131;
  assign n21133 = n6025 & n21132;
  assign n21134 = n6021 & n21133;
  assign n21135 = pi146 & ~n501;
  assign n21136 = n5713 & n21135;
  assign n21137 = n6138 & n21136;
  assign n21138 = n6147 & n21137;
  assign n21139 = ~n1172 & n21138;
  assign n21140 = ~n996 & n21139;
  assign n21141 = ~n2306 & n21140;
  assign n21142 = n3819 & n21141;
  assign n21143 = n3821 & n21142;
  assign n21144 = n6183 & n21143;
  assign n21145 = n19897 & n21144;
  assign n21146 = ~n6137 & n21145;
  assign n21147 = n6193 & n21146;
  assign n21148 = n6134 & n21147;
  assign n21149 = ~n21134 & ~n21148;
  assign n21150 = n21130 & n21149;
  assign n21151 = pi122 & ~n5598;
  assign n21152 = n6068 & n21151;
  assign n21153 = n6066 & n21152;
  assign n21154 = n6076 & n21153;
  assign n21155 = n6038 & n21154;
  assign n21156 = ~n6035 & n21155;
  assign n21157 = ~n5808 & n21156;
  assign n21158 = ~n5923 & n21157;
  assign n21159 = n6054 & n21158;
  assign n21160 = n6034 & n21159;
  assign n21161 = pi106 & ~n4677;
  assign n21162 = n4737 & n21161;
  assign n21163 = n4491 & n21162;
  assign n21164 = n4891 & n21163;
  assign n21165 = n5986 & n21164;
  assign n21166 = ~n5985 & n21165;
  assign n21167 = ~n4817 & n21166;
  assign n21168 = ~n4902 & n21167;
  assign n21169 = ~n5923 & n21168;
  assign n21170 = n5999 & n21169;
  assign n21171 = n5984 & n21170;
  assign n21172 = ~n21160 & ~n21171;
  assign n21173 = n5948 & n20147;
  assign n21174 = n5925 & n21173;
  assign n21175 = ~n5924 & n21174;
  assign n21176 = ~n3940 & n21175;
  assign n21177 = ~n4001 & n21176;
  assign n21178 = ~n5043 & n21177;
  assign n21179 = ~n5923 & n21178;
  assign n21180 = n5941 & n21179;
  assign n21181 = n5922 & n21180;
  assign n21182 = pi130 & ~n5769;
  assign n21183 = ~n5923 & n21182;
  assign n21184 = ~n5958 & n21183;
  assign n21185 = n6112 & n21184;
  assign n21186 = n6095 & n21185;
  assign n21187 = ~n21181 & ~n21186;
  assign n21188 = n21172 & n21187;
  assign n21189 = n21150 & n21188;
  assign po075 = ~n21108 | ~n21189;
  assign n21191 = n5897 & n20339;
  assign n21192 = n5771 & n21191;
  assign n21193 = ~n5770 & n21192;
  assign n21194 = ~n3066 & n21193;
  assign n21195 = ~n3983 & n21194;
  assign n21196 = ~n4003 & n21195;
  assign n21197 = ~n4024 & n21196;
  assign n21198 = ~n4999 & n21197;
  assign n21199 = ~n5751 & n21198;
  assign n21200 = n5825 & n21199;
  assign n21201 = n5750 & n21200;
  assign n21202 = n5837 & n18618;
  assign n21203 = n5839 & n21202;
  assign n21204 = n5836 & n21203;
  assign n21205 = ~n5834 & n21204;
  assign n21206 = ~n2242 & n21205;
  assign n21207 = ~n3095 & n21206;
  assign n21208 = ~n3997 & n21207;
  assign n21209 = ~n4003 & n21208;
  assign n21210 = ~n4837 & n21209;
  assign n21211 = ~n5822 & n21210;
  assign n21212 = ~n5833 & n21211;
  assign n21213 = n5856 & n21212;
  assign n21214 = n5832 & n21213;
  assign n21215 = pi043 & ~n1144;
  assign n21216 = ~n1115 & n21215;
  assign n21217 = n1056 & n21216;
  assign n21218 = ~n1208 & n21217;
  assign n21219 = n4920 & n21218;
  assign n21220 = n5873 & n21219;
  assign n21221 = n4932 & n21220;
  assign n21222 = ~n5865 & n21221;
  assign n21223 = ~n1372 & n21222;
  assign n21224 = ~n2243 & n21223;
  assign n21225 = ~n3104 & n21224;
  assign n21226 = ~n3971 & n21225;
  assign n21227 = ~n4003 & n21226;
  assign n21228 = ~n4872 & n21227;
  assign n21229 = ~n5801 & n21228;
  assign n21230 = ~n5864 & n21229;
  assign n21231 = n5891 & n21230;
  assign n21232 = n5863 & n21231;
  assign n21233 = ~n21214 & ~n21232;
  assign n21234 = ~n21201 & n21233;
  assign n21235 = ~n5058 & n20335;
  assign n21236 = ~n5923 & n21235;
  assign n21237 = n5966 & n21236;
  assign n21238 = ~n5911 & n20304;
  assign n21239 = ~n5909 & n21238;
  assign n21240 = n5916 & n21239;
  assign n21241 = pi139 & ~n501;
  assign n21242 = n6687 & n21241;
  assign n21243 = n6685 & n21242;
  assign n21244 = n6692 & n21243;
  assign n21245 = n6683 & n21244;
  assign n21246 = ~n1172 & n21245;
  assign n21247 = ~n1054 & n21246;
  assign n21248 = ~n996 & n21247;
  assign n21249 = n6698 & n21248;
  assign n21250 = n6677 & n21249;
  assign n21251 = n6707 & n21250;
  assign n21252 = n6711 & n21251;
  assign n21253 = n6676 & n21252;
  assign n21254 = n6284 & n21253;
  assign n21255 = ~n21240 & ~n21254;
  assign n21256 = ~n21237 & n21255;
  assign n21257 = ~n4881 & n20319;
  assign n21258 = ~n5923 & n21257;
  assign n21259 = n6025 & n21258;
  assign n21260 = n6021 & n21259;
  assign n21261 = pi147 & ~n501;
  assign n21262 = n5713 & n21261;
  assign n21263 = n6138 & n21262;
  assign n21264 = n6147 & n21263;
  assign n21265 = ~n1172 & n21264;
  assign n21266 = ~n996 & n21265;
  assign n21267 = ~n2306 & n21266;
  assign n21268 = n3819 & n21267;
  assign n21269 = n3821 & n21268;
  assign n21270 = n6183 & n21269;
  assign n21271 = n19897 & n21270;
  assign n21272 = ~n6137 & n21271;
  assign n21273 = n6193 & n21272;
  assign n21274 = n6134 & n21273;
  assign n21275 = ~n21260 & ~n21274;
  assign n21276 = n21256 & n21275;
  assign n21277 = pi123 & ~n5598;
  assign n21278 = n6068 & n21277;
  assign n21279 = n6066 & n21278;
  assign n21280 = n6076 & n21279;
  assign n21281 = n6038 & n21280;
  assign n21282 = ~n6035 & n21281;
  assign n21283 = ~n5808 & n21282;
  assign n21284 = ~n5923 & n21283;
  assign n21285 = n6054 & n21284;
  assign n21286 = n6034 & n21285;
  assign n21287 = pi107 & ~n4677;
  assign n21288 = n4737 & n21287;
  assign n21289 = n4491 & n21288;
  assign n21290 = n4891 & n21289;
  assign n21291 = n5986 & n21290;
  assign n21292 = ~n5985 & n21291;
  assign n21293 = ~n4817 & n21292;
  assign n21294 = ~n4902 & n21293;
  assign n21295 = ~n5923 & n21294;
  assign n21296 = n5999 & n21295;
  assign n21297 = n5984 & n21296;
  assign n21298 = ~n21286 & ~n21297;
  assign n21299 = n5948 & n20277;
  assign n21300 = n5925 & n21299;
  assign n21301 = ~n5924 & n21300;
  assign n21302 = ~n3940 & n21301;
  assign n21303 = ~n4001 & n21302;
  assign n21304 = ~n5043 & n21303;
  assign n21305 = ~n5923 & n21304;
  assign n21306 = n5941 & n21305;
  assign n21307 = n5922 & n21306;
  assign n21308 = pi131 & ~n5769;
  assign n21309 = ~n5923 & n21308;
  assign n21310 = ~n5958 & n21309;
  assign n21311 = n6112 & n21310;
  assign n21312 = n6095 & n21311;
  assign n21313 = ~n21307 & ~n21312;
  assign n21314 = n21298 & n21313;
  assign n21315 = n21276 & n21314;
  assign po076 = ~n21234 | ~n21315;
  assign n21317 = n5897 & n20443;
  assign n21318 = n5771 & n21317;
  assign n21319 = ~n5770 & n21318;
  assign n21320 = ~n3066 & n21319;
  assign n21321 = ~n3983 & n21320;
  assign n21322 = ~n4003 & n21321;
  assign n21323 = ~n4024 & n21322;
  assign n21324 = ~n4999 & n21323;
  assign n21325 = ~n5751 & n21324;
  assign n21326 = n5825 & n21325;
  assign n21327 = n5750 & n21326;
  assign n21328 = n5837 & n18656;
  assign n21329 = n5839 & n21328;
  assign n21330 = n5836 & n21329;
  assign n21331 = ~n5834 & n21330;
  assign n21332 = ~n2242 & n21331;
  assign n21333 = ~n3095 & n21332;
  assign n21334 = ~n3997 & n21333;
  assign n21335 = ~n4003 & n21334;
  assign n21336 = ~n4837 & n21335;
  assign n21337 = ~n5822 & n21336;
  assign n21338 = ~n5833 & n21337;
  assign n21339 = n5856 & n21338;
  assign n21340 = n5832 & n21339;
  assign n21341 = pi044 & ~n1144;
  assign n21342 = ~n1115 & n21341;
  assign n21343 = n1056 & n21342;
  assign n21344 = ~n1208 & n21343;
  assign n21345 = n4920 & n21344;
  assign n21346 = n5873 & n21345;
  assign n21347 = n4932 & n21346;
  assign n21348 = ~n5865 & n21347;
  assign n21349 = ~n1372 & n21348;
  assign n21350 = ~n2243 & n21349;
  assign n21351 = ~n3104 & n21350;
  assign n21352 = ~n3971 & n21351;
  assign n21353 = ~n4003 & n21352;
  assign n21354 = ~n4872 & n21353;
  assign n21355 = ~n5801 & n21354;
  assign n21356 = ~n5864 & n21355;
  assign n21357 = n5891 & n21356;
  assign n21358 = n5863 & n21357;
  assign n21359 = ~n21340 & ~n21358;
  assign n21360 = ~n21327 & n21359;
  assign n21361 = ~n5058 & n20439;
  assign n21362 = ~n5923 & n21361;
  assign n21363 = n5966 & n21362;
  assign n21364 = ~n5911 & n20408;
  assign n21365 = ~n5909 & n21364;
  assign n21366 = n5916 & n21365;
  assign n21367 = pi140 & ~n501;
  assign n21368 = n6687 & n21367;
  assign n21369 = n6685 & n21368;
  assign n21370 = n6692 & n21369;
  assign n21371 = n6683 & n21370;
  assign n21372 = ~n1172 & n21371;
  assign n21373 = ~n1054 & n21372;
  assign n21374 = ~n996 & n21373;
  assign n21375 = n6698 & n21374;
  assign n21376 = n6677 & n21375;
  assign n21377 = n6707 & n21376;
  assign n21378 = n6711 & n21377;
  assign n21379 = n6676 & n21378;
  assign n21380 = n6284 & n21379;
  assign n21381 = ~n21366 & ~n21380;
  assign n21382 = ~n21363 & n21381;
  assign n21383 = ~n4881 & n20423;
  assign n21384 = ~n5923 & n21383;
  assign n21385 = n6025 & n21384;
  assign n21386 = n6021 & n21385;
  assign n21387 = pi148 & ~n501;
  assign n21388 = n5713 & n21387;
  assign n21389 = n6138 & n21388;
  assign n21390 = n6147 & n21389;
  assign n21391 = ~n1172 & n21390;
  assign n21392 = ~n996 & n21391;
  assign n21393 = ~n2306 & n21392;
  assign n21394 = n3819 & n21393;
  assign n21395 = n3821 & n21394;
  assign n21396 = n6183 & n21395;
  assign n21397 = n19897 & n21396;
  assign n21398 = ~n6137 & n21397;
  assign n21399 = n6193 & n21398;
  assign n21400 = n6134 & n21399;
  assign n21401 = ~n21386 & ~n21400;
  assign n21402 = n21382 & n21401;
  assign n21403 = pi124 & ~n5598;
  assign n21404 = n6068 & n21403;
  assign n21405 = n6066 & n21404;
  assign n21406 = n6076 & n21405;
  assign n21407 = n6038 & n21406;
  assign n21408 = ~n6035 & n21407;
  assign n21409 = ~n5808 & n21408;
  assign n21410 = ~n5923 & n21409;
  assign n21411 = n6054 & n21410;
  assign n21412 = n6034 & n21411;
  assign n21413 = pi108 & ~n4677;
  assign n21414 = n4737 & n21413;
  assign n21415 = n4491 & n21414;
  assign n21416 = n4891 & n21415;
  assign n21417 = n5986 & n21416;
  assign n21418 = ~n5985 & n21417;
  assign n21419 = ~n4817 & n21418;
  assign n21420 = ~n4902 & n21419;
  assign n21421 = ~n5923 & n21420;
  assign n21422 = n5999 & n21421;
  assign n21423 = n5984 & n21422;
  assign n21424 = ~n21412 & ~n21423;
  assign n21425 = n5948 & n20381;
  assign n21426 = n5925 & n21425;
  assign n21427 = ~n5924 & n21426;
  assign n21428 = ~n3940 & n21427;
  assign n21429 = ~n4001 & n21428;
  assign n21430 = ~n5043 & n21429;
  assign n21431 = ~n5923 & n21430;
  assign n21432 = n5941 & n21431;
  assign n21433 = n5922 & n21432;
  assign n21434 = pi132 & ~n5769;
  assign n21435 = ~n5923 & n21434;
  assign n21436 = ~n5958 & n21435;
  assign n21437 = n6112 & n21436;
  assign n21438 = n6095 & n21437;
  assign n21439 = ~n21433 & ~n21438;
  assign n21440 = n21424 & n21439;
  assign n21441 = n21402 & n21440;
  assign po077 = ~n21360 | ~n21441;
  assign n21443 = n5897 & n20547;
  assign n21444 = n5771 & n21443;
  assign n21445 = ~n5770 & n21444;
  assign n21446 = ~n3066 & n21445;
  assign n21447 = ~n3983 & n21446;
  assign n21448 = ~n4003 & n21447;
  assign n21449 = ~n4024 & n21448;
  assign n21450 = ~n4999 & n21449;
  assign n21451 = ~n5751 & n21450;
  assign n21452 = n5825 & n21451;
  assign n21453 = n5750 & n21452;
  assign n21454 = n5837 & n18694;
  assign n21455 = n5839 & n21454;
  assign n21456 = n5836 & n21455;
  assign n21457 = ~n5834 & n21456;
  assign n21458 = ~n2242 & n21457;
  assign n21459 = ~n3095 & n21458;
  assign n21460 = ~n3997 & n21459;
  assign n21461 = ~n4003 & n21460;
  assign n21462 = ~n4837 & n21461;
  assign n21463 = ~n5822 & n21462;
  assign n21464 = ~n5833 & n21463;
  assign n21465 = n5856 & n21464;
  assign n21466 = n5832 & n21465;
  assign n21467 = pi045 & ~n1144;
  assign n21468 = ~n1115 & n21467;
  assign n21469 = n1056 & n21468;
  assign n21470 = ~n1208 & n21469;
  assign n21471 = n4920 & n21470;
  assign n21472 = n5873 & n21471;
  assign n21473 = n4932 & n21472;
  assign n21474 = ~n5865 & n21473;
  assign n21475 = ~n1372 & n21474;
  assign n21476 = ~n2243 & n21475;
  assign n21477 = ~n3104 & n21476;
  assign n21478 = ~n3971 & n21477;
  assign n21479 = ~n4003 & n21478;
  assign n21480 = ~n4872 & n21479;
  assign n21481 = ~n5801 & n21480;
  assign n21482 = ~n5864 & n21481;
  assign n21483 = n5891 & n21482;
  assign n21484 = n5863 & n21483;
  assign n21485 = ~n21466 & ~n21484;
  assign n21486 = ~n21453 & n21485;
  assign n21487 = ~n5058 & n20543;
  assign n21488 = ~n5923 & n21487;
  assign n21489 = n5966 & n21488;
  assign n21490 = ~n5911 & n20512;
  assign n21491 = ~n5909 & n21490;
  assign n21492 = n5916 & n21491;
  assign n21493 = pi141 & ~n501;
  assign n21494 = n6687 & n21493;
  assign n21495 = n6685 & n21494;
  assign n21496 = n6692 & n21495;
  assign n21497 = n6683 & n21496;
  assign n21498 = ~n1172 & n21497;
  assign n21499 = ~n1054 & n21498;
  assign n21500 = ~n996 & n21499;
  assign n21501 = n6698 & n21500;
  assign n21502 = n6677 & n21501;
  assign n21503 = n6707 & n21502;
  assign n21504 = n6711 & n21503;
  assign n21505 = n6676 & n21504;
  assign n21506 = n6284 & n21505;
  assign n21507 = ~n21492 & ~n21506;
  assign n21508 = ~n21489 & n21507;
  assign n21509 = ~n4881 & n20527;
  assign n21510 = ~n5923 & n21509;
  assign n21511 = n6025 & n21510;
  assign n21512 = n6021 & n21511;
  assign n21513 = pi149 & ~n501;
  assign n21514 = n5713 & n21513;
  assign n21515 = n6138 & n21514;
  assign n21516 = n6147 & n21515;
  assign n21517 = ~n1172 & n21516;
  assign n21518 = ~n996 & n21517;
  assign n21519 = ~n2306 & n21518;
  assign n21520 = n3819 & n21519;
  assign n21521 = n3821 & n21520;
  assign n21522 = n6183 & n21521;
  assign n21523 = n19897 & n21522;
  assign n21524 = ~n6137 & n21523;
  assign n21525 = n6193 & n21524;
  assign n21526 = n6134 & n21525;
  assign n21527 = ~n21512 & ~n21526;
  assign n21528 = n21508 & n21527;
  assign n21529 = pi125 & ~n5598;
  assign n21530 = n6068 & n21529;
  assign n21531 = n6066 & n21530;
  assign n21532 = n6076 & n21531;
  assign n21533 = n6038 & n21532;
  assign n21534 = ~n6035 & n21533;
  assign n21535 = ~n5808 & n21534;
  assign n21536 = ~n5923 & n21535;
  assign n21537 = n6054 & n21536;
  assign n21538 = n6034 & n21537;
  assign n21539 = pi109 & ~n4677;
  assign n21540 = n4737 & n21539;
  assign n21541 = n4491 & n21540;
  assign n21542 = n4891 & n21541;
  assign n21543 = n5986 & n21542;
  assign n21544 = ~n5985 & n21543;
  assign n21545 = ~n4817 & n21544;
  assign n21546 = ~n4902 & n21545;
  assign n21547 = ~n5923 & n21546;
  assign n21548 = n5999 & n21547;
  assign n21549 = n5984 & n21548;
  assign n21550 = ~n21538 & ~n21549;
  assign n21551 = n5948 & n20485;
  assign n21552 = n5925 & n21551;
  assign n21553 = ~n5924 & n21552;
  assign n21554 = ~n3940 & n21553;
  assign n21555 = ~n4001 & n21554;
  assign n21556 = ~n5043 & n21555;
  assign n21557 = ~n5923 & n21556;
  assign n21558 = n5941 & n21557;
  assign n21559 = n5922 & n21558;
  assign n21560 = pi133 & ~n5769;
  assign n21561 = ~n5923 & n21560;
  assign n21562 = ~n5958 & n21561;
  assign n21563 = n6112 & n21562;
  assign n21564 = n6095 & n21563;
  assign n21565 = ~n21559 & ~n21564;
  assign n21566 = n21550 & n21565;
  assign n21567 = n21528 & n21566;
  assign po078 = ~n21486 | ~n21567;
  assign n21569 = n5897 & n20651;
  assign n21570 = n5771 & n21569;
  assign n21571 = ~n5770 & n21570;
  assign n21572 = ~n3066 & n21571;
  assign n21573 = ~n3983 & n21572;
  assign n21574 = ~n4003 & n21573;
  assign n21575 = ~n4024 & n21574;
  assign n21576 = ~n4999 & n21575;
  assign n21577 = ~n5751 & n21576;
  assign n21578 = n5825 & n21577;
  assign n21579 = n5750 & n21578;
  assign n21580 = n5837 & n18732;
  assign n21581 = n5839 & n21580;
  assign n21582 = n5836 & n21581;
  assign n21583 = ~n5834 & n21582;
  assign n21584 = ~n2242 & n21583;
  assign n21585 = ~n3095 & n21584;
  assign n21586 = ~n3997 & n21585;
  assign n21587 = ~n4003 & n21586;
  assign n21588 = ~n4837 & n21587;
  assign n21589 = ~n5822 & n21588;
  assign n21590 = ~n5833 & n21589;
  assign n21591 = n5856 & n21590;
  assign n21592 = n5832 & n21591;
  assign n21593 = pi046 & ~n1144;
  assign n21594 = ~n1115 & n21593;
  assign n21595 = n1056 & n21594;
  assign n21596 = ~n1208 & n21595;
  assign n21597 = n4920 & n21596;
  assign n21598 = n5873 & n21597;
  assign n21599 = n4932 & n21598;
  assign n21600 = ~n5865 & n21599;
  assign n21601 = ~n1372 & n21600;
  assign n21602 = ~n2243 & n21601;
  assign n21603 = ~n3104 & n21602;
  assign n21604 = ~n3971 & n21603;
  assign n21605 = ~n4003 & n21604;
  assign n21606 = ~n4872 & n21605;
  assign n21607 = ~n5801 & n21606;
  assign n21608 = ~n5864 & n21607;
  assign n21609 = n5891 & n21608;
  assign n21610 = n5863 & n21609;
  assign n21611 = ~n21592 & ~n21610;
  assign n21612 = ~n21579 & n21611;
  assign n21613 = ~n5058 & n20647;
  assign n21614 = ~n5923 & n21613;
  assign n21615 = n5966 & n21614;
  assign n21616 = ~n5911 & n20616;
  assign n21617 = ~n5909 & n21616;
  assign n21618 = n5916 & n21617;
  assign n21619 = pi142 & ~n501;
  assign n21620 = n6687 & n21619;
  assign n21621 = n6685 & n21620;
  assign n21622 = n6692 & n21621;
  assign n21623 = n6683 & n21622;
  assign n21624 = ~n1172 & n21623;
  assign n21625 = ~n1054 & n21624;
  assign n21626 = ~n996 & n21625;
  assign n21627 = n6698 & n21626;
  assign n21628 = n6677 & n21627;
  assign n21629 = n6707 & n21628;
  assign n21630 = n6711 & n21629;
  assign n21631 = n6676 & n21630;
  assign n21632 = n6284 & n21631;
  assign n21633 = ~n21618 & ~n21632;
  assign n21634 = ~n21615 & n21633;
  assign n21635 = ~n4881 & n20631;
  assign n21636 = ~n5923 & n21635;
  assign n21637 = n6025 & n21636;
  assign n21638 = n6021 & n21637;
  assign n21639 = pi150 & ~n501;
  assign n21640 = n5713 & n21639;
  assign n21641 = n6138 & n21640;
  assign n21642 = n6147 & n21641;
  assign n21643 = ~n1172 & n21642;
  assign n21644 = ~n996 & n21643;
  assign n21645 = ~n2306 & n21644;
  assign n21646 = n3819 & n21645;
  assign n21647 = n3821 & n21646;
  assign n21648 = n6183 & n21647;
  assign n21649 = n19897 & n21648;
  assign n21650 = ~n6137 & n21649;
  assign n21651 = n6193 & n21650;
  assign n21652 = n6134 & n21651;
  assign n21653 = ~n21638 & ~n21652;
  assign n21654 = n21634 & n21653;
  assign n21655 = pi126 & ~n5598;
  assign n21656 = n6068 & n21655;
  assign n21657 = n6066 & n21656;
  assign n21658 = n6076 & n21657;
  assign n21659 = n6038 & n21658;
  assign n21660 = ~n6035 & n21659;
  assign n21661 = ~n5808 & n21660;
  assign n21662 = ~n5923 & n21661;
  assign n21663 = n6054 & n21662;
  assign n21664 = n6034 & n21663;
  assign n21665 = pi110 & ~n4677;
  assign n21666 = n4737 & n21665;
  assign n21667 = n4491 & n21666;
  assign n21668 = n4891 & n21667;
  assign n21669 = n5986 & n21668;
  assign n21670 = ~n5985 & n21669;
  assign n21671 = ~n4817 & n21670;
  assign n21672 = ~n4902 & n21671;
  assign n21673 = ~n5923 & n21672;
  assign n21674 = n5999 & n21673;
  assign n21675 = n5984 & n21674;
  assign n21676 = ~n21664 & ~n21675;
  assign n21677 = n5948 & n20589;
  assign n21678 = n5925 & n21677;
  assign n21679 = ~n5924 & n21678;
  assign n21680 = ~n3940 & n21679;
  assign n21681 = ~n4001 & n21680;
  assign n21682 = ~n5043 & n21681;
  assign n21683 = ~n5923 & n21682;
  assign n21684 = n5941 & n21683;
  assign n21685 = n5922 & n21684;
  assign n21686 = pi134 & ~n5769;
  assign n21687 = ~n5923 & n21686;
  assign n21688 = ~n5958 & n21687;
  assign n21689 = n6112 & n21688;
  assign n21690 = n6095 & n21689;
  assign n21691 = ~n21685 & ~n21690;
  assign n21692 = n21676 & n21691;
  assign n21693 = n21654 & n21692;
  assign po079 = ~n21612 | ~n21693;
  assign n21695 = pi135 & ~n6432;
  assign n21696 = n7170 & n21695;
  assign n21697 = n7178 & n21696;
  assign n21698 = n6284 & n21697;
  assign n21699 = ~n6784 & n21698;
  assign n21700 = ~n6931 & n21699;
  assign n21701 = ~n6959 & n21700;
  assign n21702 = n7142 & n21701;
  assign n21703 = n7156 & n21702;
  assign n21704 = n7132 & n21703;
  assign n21705 = pi143 & ~n7193;
  assign n21706 = ~n6754 & n21705;
  assign n21707 = ~n6931 & n21706;
  assign n21708 = n7054 & n21707;
  assign n21709 = n7202 & n21708;
  assign n21710 = n7192 & n21709;
  assign n21711 = ~n2543 & n20790;
  assign n21712 = n5772 & n21711;
  assign n21713 = ~n2842 & n3850;
  assign n21714 = n5775 & n21713;
  assign n21715 = n21712 & n21714;
  assign n21716 = n6875 & n21715;
  assign n21717 = ~n6874 & n21716;
  assign n21718 = ~n3066 & n21717;
  assign n21719 = ~n3983 & n21718;
  assign n21720 = ~n4003 & n21719;
  assign n21721 = ~n4024 & n21720;
  assign n21722 = ~n4999 & n21721;
  assign n21723 = ~n6873 & n21722;
  assign n21724 = ~n5827 & n21723;
  assign n21725 = ~n6872 & n21724;
  assign n21726 = n6890 & n21725;
  assign n21727 = n6871 & n21726;
  assign n21728 = n6866 & n21727;
  assign n21729 = ~n21710 & ~n21728;
  assign n21730 = ~n21704 & n21729;
  assign n21731 = n7030 & n20696;
  assign n21732 = n7034 & n21731;
  assign n21733 = n6998 & n21732;
  assign n21734 = ~n6997 & n21733;
  assign n21735 = ~n4817 & n21734;
  assign n21736 = ~n4902 & n21735;
  assign n21737 = ~n6931 & n21736;
  assign n21738 = ~n6001 & n21737;
  assign n21739 = ~n6996 & n21738;
  assign n21740 = n7011 & n21739;
  assign n21741 = n6995 & n21740;
  assign n21742 = n6991 & n21741;
  assign n21743 = ~n1026 & n20752;
  assign n21744 = n6787 & n21743;
  assign n21745 = n1239 & n21744;
  assign n21746 = ~n1270 & n21745;
  assign n21747 = n844 & n21746;
  assign n21748 = ~n1372 & n21747;
  assign n21749 = ~n2243 & n21748;
  assign n21750 = ~n6785 & n21749;
  assign n21751 = ~n3104 & n21750;
  assign n21752 = ~n3971 & n21751;
  assign n21753 = ~n4003 & n21752;
  assign n21754 = ~n4872 & n21753;
  assign n21755 = ~n5801 & n21754;
  assign n21756 = ~n6761 & n21755;
  assign n21757 = ~n6760 & n21756;
  assign n21758 = ~n6759 & n21757;
  assign n21759 = n6822 & n21758;
  assign n21760 = n6758 & n21759;
  assign n21761 = n6722 & n21760;
  assign n21762 = ~n21742 & ~n21761;
  assign n21763 = n3800 & n20682;
  assign n21764 = n3681 & n5947;
  assign n21765 = n21763 & n21764;
  assign n21766 = n6934 & n21765;
  assign n21767 = ~n6932 & n21766;
  assign n21768 = ~n3940 & n21767;
  assign n21769 = ~n4001 & n21768;
  assign n21770 = ~n5043 & n21769;
  assign n21771 = ~n6931 & n21770;
  assign n21772 = ~n5943 & n21771;
  assign n21773 = ~n6930 & n21772;
  assign n21774 = n6948 & n21773;
  assign n21775 = n6929 & n21774;
  assign n21776 = n6924 & n21775;
  assign n21777 = n7096 & n20774;
  assign n21778 = n6074 & n20777;
  assign n21779 = n7099 & n21778;
  assign n21780 = n6036 & n21779;
  assign n21781 = n21777 & n21780;
  assign n21782 = ~n7057 & n21781;
  assign n21783 = ~n5808 & n21782;
  assign n21784 = ~n6931 & n21783;
  assign n21785 = ~n6056 & n21784;
  assign n21786 = ~n7056 & n21785;
  assign n21787 = n7070 & n21786;
  assign n21788 = n7055 & n21787;
  assign n21789 = n7052 & n21788;
  assign n21790 = ~n21776 & ~n21789;
  assign n21791 = n21762 & n21790;
  assign n21792 = ~n5967 & n20742;
  assign n21793 = ~n6931 & n21792;
  assign n21794 = ~n6958 & n21793;
  assign n21795 = n6966 & n21794;
  assign n21796 = ~n6027 & n20745;
  assign n21797 = ~n6931 & n21796;
  assign n21798 = ~n6959 & n21797;
  assign n21799 = n7027 & n21798;
  assign n21800 = n7021 & n21799;
  assign n21801 = ~n6931 & n20804;
  assign n21802 = ~n6114 & n21801;
  assign n21803 = n7054 & n21802;
  assign n21804 = n7093 & n21803;
  assign n21805 = n7087 & n21804;
  assign n21806 = ~n21800 & ~n21805;
  assign n21807 = ~n21795 & n21806;
  assign n21808 = n5835 & n18802;
  assign n21809 = n6843 & n21808;
  assign n21810 = ~n6838 & n21809;
  assign n21811 = ~n2242 & n21810;
  assign n21812 = ~n3095 & n21811;
  assign n21813 = ~n3997 & n21812;
  assign n21814 = ~n4003 & n21813;
  assign n21815 = ~n4837 & n21814;
  assign n21816 = ~n5822 & n21815;
  assign n21817 = ~n6837 & n21816;
  assign n21818 = ~n6820 & n21817;
  assign n21819 = ~n6836 & n21818;
  assign n21820 = n6857 & n21819;
  assign n21821 = n6835 & n21820;
  assign n21822 = n6830 & n21821;
  assign n21823 = pi159 & ~n501;
  assign n21824 = n5713 & n21823;
  assign n21825 = n6138 & n21824;
  assign n21826 = n7244 & n21825;
  assign n21827 = ~n1172 & n21826;
  assign n21828 = ~n996 & n21827;
  assign n21829 = ~n2306 & n21828;
  assign n21830 = ~n500 & n21829;
  assign n21831 = n6677 & n21830;
  assign n21832 = n7280 & n21831;
  assign n21833 = n7284 & n21832;
  assign n21834 = ~n7236 & n21833;
  assign n21835 = ~n6137 & n21834;
  assign n21836 = n6193 & n21835;
  assign n21837 = n6134 & n21836;
  assign n21838 = ~n7235 & n21837;
  assign n21839 = n7296 & n21838;
  assign n21840 = n7231 & n21839;
  assign n21841 = ~n5917 & n20723;
  assign n21842 = ~n6911 & n21841;
  assign n21843 = n6916 & n21842;
  assign n21844 = ~n2812 & ~n3254;
  assign n21845 = n7598 & n21844;
  assign n21846 = n3819 & n18099;
  assign n21847 = n21845 & n21846;
  assign n21848 = n7606 & n21847;
  assign n21849 = pi151 & ~n501;
  assign n21850 = n7621 & n21849;
  assign n21851 = n7625 & n21850;
  assign n21852 = n7618 & n21851;
  assign n21853 = ~n1172 & n21852;
  assign n21854 = ~n1143 & n21853;
  assign n21855 = ~n996 & n21854;
  assign n21856 = ~n2306 & n21855;
  assign n21857 = ~n500 & n21856;
  assign n21858 = n2316 & n21857;
  assign n21859 = n7608 & n21858;
  assign n21860 = n7757 & n21859;
  assign n21861 = n21848 & n21860;
  assign n21862 = n7597 & n21861;
  assign n21863 = ~n6137 & n21862;
  assign n21864 = n6193 & n21863;
  assign n21865 = n6134 & n21864;
  assign n21866 = ~n21843 & ~n21865;
  assign n21867 = ~n21840 & n21866;
  assign n21868 = ~n21822 & n21867;
  assign n21869 = n21807 & n21868;
  assign n21870 = n21791 & n21869;
  assign po080 = ~n21730 | ~n21870;
  assign n21872 = n7096 & n20899;
  assign n21873 = n7100 & n21872;
  assign n21874 = n7058 & n21873;
  assign n21875 = ~n7057 & n21874;
  assign n21876 = ~n5808 & n21875;
  assign n21877 = ~n6931 & n21876;
  assign n21878 = ~n6056 & n21877;
  assign n21879 = ~n7056 & n21878;
  assign n21880 = n7070 & n21879;
  assign n21881 = n7055 & n21880;
  assign n21882 = n7052 & n21881;
  assign n21883 = pi072 & ~n2543;
  assign n21884 = n5772 & n21883;
  assign n21885 = n5776 & n21884;
  assign n21886 = n6875 & n21885;
  assign n21887 = ~n6874 & n21886;
  assign n21888 = ~n3066 & n21887;
  assign n21889 = ~n3983 & n21888;
  assign n21890 = ~n4003 & n21889;
  assign n21891 = ~n4024 & n21890;
  assign n21892 = ~n4999 & n21891;
  assign n21893 = ~n6873 & n21892;
  assign n21894 = ~n5827 & n21893;
  assign n21895 = ~n6872 & n21894;
  assign n21896 = n6890 & n21895;
  assign n21897 = n6871 & n21896;
  assign n21898 = n6866 & n21897;
  assign n21899 = pi144 & ~n7193;
  assign n21900 = ~n6754 & n21899;
  assign n21901 = ~n6931 & n21900;
  assign n21902 = n7054 & n21901;
  assign n21903 = n7202 & n21902;
  assign n21904 = n7192 & n21903;
  assign n21905 = ~n21898 & ~n21904;
  assign n21906 = ~n21882 & n21905;
  assign n21907 = n5835 & n18861;
  assign n21908 = n6843 & n21907;
  assign n21909 = ~n6838 & n21908;
  assign n21910 = ~n2242 & n21909;
  assign n21911 = ~n3095 & n21910;
  assign n21912 = ~n3997 & n21911;
  assign n21913 = ~n4003 & n21912;
  assign n21914 = ~n4837 & n21913;
  assign n21915 = ~n5822 & n21914;
  assign n21916 = ~n6837 & n21915;
  assign n21917 = ~n6820 & n21916;
  assign n21918 = ~n6836 & n21917;
  assign n21919 = n6857 & n21918;
  assign n21920 = n6835 & n21919;
  assign n21921 = n6830 & n21920;
  assign n21922 = n3800 & n19386;
  assign n21923 = n5927 & n21922;
  assign n21924 = n6934 & n21923;
  assign n21925 = ~n6932 & n21924;
  assign n21926 = ~n3940 & n21925;
  assign n21927 = ~n4001 & n21926;
  assign n21928 = ~n5043 & n21927;
  assign n21929 = ~n6931 & n21928;
  assign n21930 = ~n5943 & n21929;
  assign n21931 = ~n6930 & n21930;
  assign n21932 = n6948 & n21931;
  assign n21933 = n6929 & n21932;
  assign n21934 = n6924 & n21933;
  assign n21935 = ~n21921 & ~n21934;
  assign n21936 = n7030 & n20844;
  assign n21937 = n7034 & n21936;
  assign n21938 = n6998 & n21937;
  assign n21939 = ~n6997 & n21938;
  assign n21940 = ~n4817 & n21939;
  assign n21941 = ~n4902 & n21940;
  assign n21942 = ~n6931 & n21941;
  assign n21943 = ~n6001 & n21942;
  assign n21944 = ~n6996 & n21943;
  assign n21945 = n7011 & n21944;
  assign n21946 = n6995 & n21945;
  assign n21947 = n6991 & n21946;
  assign n21948 = pi136 & ~n6432;
  assign n21949 = n7170 & n21948;
  assign n21950 = n7178 & n21949;
  assign n21951 = n6284 & n21950;
  assign n21952 = ~n6784 & n21951;
  assign n21953 = ~n6931 & n21952;
  assign n21954 = ~n6959 & n21953;
  assign n21955 = n7142 & n21954;
  assign n21956 = n7156 & n21955;
  assign n21957 = n7132 & n21956;
  assign n21958 = ~n21947 & ~n21957;
  assign n21959 = n21935 & n21958;
  assign n21960 = ~n6931 & n20919;
  assign n21961 = ~n6114 & n21960;
  assign n21962 = n7054 & n21961;
  assign n21963 = n7093 & n21962;
  assign n21964 = n7087 & n21963;
  assign n21965 = ~n6027 & n20879;
  assign n21966 = ~n6931 & n21965;
  assign n21967 = ~n6959 & n21966;
  assign n21968 = n7027 & n21967;
  assign n21969 = n7021 & n21968;
  assign n21970 = ~n5967 & n20857;
  assign n21971 = ~n6931 & n21970;
  assign n21972 = ~n6958 & n21971;
  assign n21973 = n6966 & n21972;
  assign n21974 = ~n21969 & ~n21973;
  assign n21975 = ~n21964 & n21974;
  assign n21976 = ~n1026 & n20814;
  assign n21977 = n6787 & n21976;
  assign n21978 = n1239 & n21977;
  assign n21979 = ~n1270 & n21978;
  assign n21980 = n844 & n21979;
  assign n21981 = ~n1372 & n21980;
  assign n21982 = ~n2243 & n21981;
  assign n21983 = ~n6785 & n21982;
  assign n21984 = ~n3104 & n21983;
  assign n21985 = ~n3971 & n21984;
  assign n21986 = ~n4003 & n21985;
  assign n21987 = ~n4872 & n21986;
  assign n21988 = ~n5801 & n21987;
  assign n21989 = ~n6761 & n21988;
  assign n21990 = ~n6760 & n21989;
  assign n21991 = ~n6759 & n21990;
  assign n21992 = n6822 & n21991;
  assign n21993 = n6758 & n21992;
  assign n21994 = n6722 & n21993;
  assign n21995 = pi160 & ~n501;
  assign n21996 = n5713 & n21995;
  assign n21997 = n6138 & n21996;
  assign n21998 = n7244 & n21997;
  assign n21999 = ~n1172 & n21998;
  assign n22000 = ~n996 & n21999;
  assign n22001 = ~n2306 & n22000;
  assign n22002 = ~n500 & n22001;
  assign n22003 = n6677 & n22002;
  assign n22004 = n7280 & n22003;
  assign n22005 = n7284 & n22004;
  assign n22006 = ~n7236 & n22005;
  assign n22007 = ~n6137 & n22006;
  assign n22008 = n6193 & n22007;
  assign n22009 = n6134 & n22008;
  assign n22010 = ~n7235 & n22009;
  assign n22011 = n7296 & n22010;
  assign n22012 = n7231 & n22011;
  assign n22013 = ~n5917 & n20860;
  assign n22014 = ~n6911 & n22013;
  assign n22015 = n6916 & n22014;
  assign n22016 = pi152 & ~n501;
  assign n22017 = n7621 & n22016;
  assign n22018 = n7625 & n22017;
  assign n22019 = n7618 & n22018;
  assign n22020 = ~n1172 & n22019;
  assign n22021 = ~n1143 & n22020;
  assign n22022 = ~n996 & n22021;
  assign n22023 = ~n2306 & n22022;
  assign n22024 = ~n500 & n22023;
  assign n22025 = n2316 & n22024;
  assign n22026 = n7608 & n22025;
  assign n22027 = n7757 & n22026;
  assign n22028 = n21848 & n22027;
  assign n22029 = n7597 & n22028;
  assign n22030 = ~n6137 & n22029;
  assign n22031 = n6193 & n22030;
  assign n22032 = n6134 & n22031;
  assign n22033 = ~n22015 & ~n22032;
  assign n22034 = ~n22012 & n22033;
  assign n22035 = ~n21994 & n22034;
  assign n22036 = n21975 & n22035;
  assign n22037 = n21959 & n22036;
  assign po081 = ~n21906 | ~n22037;
  assign n22039 = pi145 & ~n7193;
  assign n22040 = ~n6754 & n22039;
  assign n22041 = ~n6931 & n22040;
  assign n22042 = n7054 & n22041;
  assign n22043 = n7202 & n22042;
  assign n22044 = n7192 & n22043;
  assign n22045 = pi137 & ~n6432;
  assign n22046 = n7170 & n22045;
  assign n22047 = n7178 & n22046;
  assign n22048 = n6284 & n22047;
  assign n22049 = ~n6784 & n22048;
  assign n22050 = ~n6931 & n22049;
  assign n22051 = ~n6959 & n22050;
  assign n22052 = n7142 & n22051;
  assign n22053 = n7156 & n22052;
  assign n22054 = n7132 & n22053;
  assign n22055 = pi073 & ~n2543;
  assign n22056 = n5772 & n22055;
  assign n22057 = n5776 & n22056;
  assign n22058 = n6875 & n22057;
  assign n22059 = ~n6874 & n22058;
  assign n22060 = ~n3066 & n22059;
  assign n22061 = ~n3983 & n22060;
  assign n22062 = ~n4003 & n22061;
  assign n22063 = ~n4024 & n22062;
  assign n22064 = ~n4999 & n22063;
  assign n22065 = ~n6873 & n22064;
  assign n22066 = ~n5827 & n22065;
  assign n22067 = ~n6872 & n22066;
  assign n22068 = n6890 & n22067;
  assign n22069 = n6871 & n22068;
  assign n22070 = n6866 & n22069;
  assign n22071 = ~n22054 & ~n22070;
  assign n22072 = ~n22044 & n22071;
  assign n22073 = n7096 & n21025;
  assign n22074 = n7100 & n22073;
  assign n22075 = n7058 & n22074;
  assign n22076 = ~n7057 & n22075;
  assign n22077 = ~n5808 & n22076;
  assign n22078 = ~n6931 & n22077;
  assign n22079 = ~n6056 & n22078;
  assign n22080 = ~n7056 & n22079;
  assign n22081 = n7070 & n22080;
  assign n22082 = n7055 & n22081;
  assign n22083 = n7052 & n22082;
  assign n22084 = n5835 & n18933;
  assign n22085 = n6843 & n22084;
  assign n22086 = ~n6838 & n22085;
  assign n22087 = ~n2242 & n22086;
  assign n22088 = ~n3095 & n22087;
  assign n22089 = ~n3997 & n22088;
  assign n22090 = ~n4003 & n22089;
  assign n22091 = ~n4837 & n22090;
  assign n22092 = ~n5822 & n22091;
  assign n22093 = ~n6837 & n22092;
  assign n22094 = ~n6820 & n22093;
  assign n22095 = ~n6836 & n22094;
  assign n22096 = n6857 & n22095;
  assign n22097 = n6835 & n22096;
  assign n22098 = n6830 & n22097;
  assign n22099 = ~n22083 & ~n22098;
  assign n22100 = ~n1026 & n20964;
  assign n22101 = n6787 & n22100;
  assign n22102 = n1239 & n22101;
  assign n22103 = ~n1270 & n22102;
  assign n22104 = n844 & n22103;
  assign n22105 = ~n1372 & n22104;
  assign n22106 = ~n2243 & n22105;
  assign n22107 = ~n6785 & n22106;
  assign n22108 = ~n3104 & n22107;
  assign n22109 = ~n3971 & n22108;
  assign n22110 = ~n4003 & n22109;
  assign n22111 = ~n4872 & n22110;
  assign n22112 = ~n5801 & n22111;
  assign n22113 = ~n6761 & n22112;
  assign n22114 = ~n6760 & n22113;
  assign n22115 = ~n6759 & n22114;
  assign n22116 = n6822 & n22115;
  assign n22117 = n6758 & n22116;
  assign n22118 = n6722 & n22117;
  assign n22119 = n7030 & n21035;
  assign n22120 = n7034 & n22119;
  assign n22121 = n6998 & n22120;
  assign n22122 = ~n6997 & n22121;
  assign n22123 = ~n4817 & n22122;
  assign n22124 = ~n4902 & n22123;
  assign n22125 = ~n6931 & n22124;
  assign n22126 = ~n6001 & n22125;
  assign n22127 = ~n6996 & n22126;
  assign n22128 = n7011 & n22127;
  assign n22129 = n6995 & n22128;
  assign n22130 = n6991 & n22129;
  assign n22131 = ~n22118 & ~n22130;
  assign n22132 = n22099 & n22131;
  assign n22133 = pi161 & ~n501;
  assign n22134 = n5713 & n22133;
  assign n22135 = n6138 & n22134;
  assign n22136 = n7244 & n22135;
  assign n22137 = ~n1172 & n22136;
  assign n22138 = ~n996 & n22137;
  assign n22139 = ~n2306 & n22138;
  assign n22140 = ~n500 & n22139;
  assign n22141 = n6677 & n22140;
  assign n22142 = n7280 & n22141;
  assign n22143 = n7284 & n22142;
  assign n22144 = ~n7236 & n22143;
  assign n22145 = ~n6137 & n22144;
  assign n22146 = n6193 & n22145;
  assign n22147 = n6134 & n22146;
  assign n22148 = ~n7235 & n22147;
  assign n22149 = n7296 & n22148;
  assign n22150 = n7231 & n22149;
  assign n22151 = ~n6027 & n21005;
  assign n22152 = ~n6931 & n22151;
  assign n22153 = ~n6959 & n22152;
  assign n22154 = n7027 & n22153;
  assign n22155 = n7021 & n22154;
  assign n22156 = ~n6931 & n21056;
  assign n22157 = ~n6114 & n22156;
  assign n22158 = n7054 & n22157;
  assign n22159 = n7093 & n22158;
  assign n22160 = n7087 & n22159;
  assign n22161 = ~n22155 & ~n22160;
  assign n22162 = ~n22150 & n22161;
  assign n22163 = n3800 & n19437;
  assign n22164 = n5927 & n22163;
  assign n22165 = n6934 & n22164;
  assign n22166 = ~n6932 & n22165;
  assign n22167 = ~n3940 & n22166;
  assign n22168 = ~n4001 & n22167;
  assign n22169 = ~n5043 & n22168;
  assign n22170 = ~n6931 & n22169;
  assign n22171 = ~n5943 & n22170;
  assign n22172 = ~n6930 & n22171;
  assign n22173 = n6948 & n22172;
  assign n22174 = n6929 & n22173;
  assign n22175 = n6924 & n22174;
  assign n22176 = ~n5967 & n20983;
  assign n22177 = ~n6931 & n22176;
  assign n22178 = ~n6958 & n22177;
  assign n22179 = n6966 & n22178;
  assign n22180 = ~n5917 & n20986;
  assign n22181 = ~n6911 & n22180;
  assign n22182 = n6916 & n22181;
  assign n22183 = pi153 & ~n501;
  assign n22184 = n7621 & n22183;
  assign n22185 = n7625 & n22184;
  assign n22186 = n7618 & n22185;
  assign n22187 = ~n1172 & n22186;
  assign n22188 = ~n1143 & n22187;
  assign n22189 = ~n996 & n22188;
  assign n22190 = ~n2306 & n22189;
  assign n22191 = ~n500 & n22190;
  assign n22192 = n2316 & n22191;
  assign n22193 = n7608 & n22192;
  assign n22194 = n7757 & n22193;
  assign n22195 = n21848 & n22194;
  assign n22196 = n7597 & n22195;
  assign n22197 = ~n6137 & n22196;
  assign n22198 = n6193 & n22197;
  assign n22199 = n6134 & n22198;
  assign n22200 = ~n22182 & ~n22199;
  assign n22201 = ~n22179 & n22200;
  assign n22202 = ~n22175 & n22201;
  assign n22203 = n22162 & n22202;
  assign n22204 = n22132 & n22203;
  assign po082 = ~n22072 | ~n22204;
  assign n22206 = ~n1026 & n21090;
  assign n22207 = n6787 & n22206;
  assign n22208 = n1239 & n22207;
  assign n22209 = ~n1270 & n22208;
  assign n22210 = n844 & n22209;
  assign n22211 = ~n1372 & n22210;
  assign n22212 = ~n2243 & n22211;
  assign n22213 = ~n6785 & n22212;
  assign n22214 = ~n3104 & n22213;
  assign n22215 = ~n3971 & n22214;
  assign n22216 = ~n4003 & n22215;
  assign n22217 = ~n4872 & n22216;
  assign n22218 = ~n5801 & n22217;
  assign n22219 = ~n6761 & n22218;
  assign n22220 = ~n6760 & n22219;
  assign n22221 = ~n6759 & n22220;
  assign n22222 = n6822 & n22221;
  assign n22223 = n6758 & n22222;
  assign n22224 = n6722 & n22223;
  assign n22225 = pi146 & ~n7193;
  assign n22226 = ~n6754 & n22225;
  assign n22227 = ~n6931 & n22226;
  assign n22228 = n7054 & n22227;
  assign n22229 = n7202 & n22228;
  assign n22230 = n7192 & n22229;
  assign n22231 = n7096 & n21151;
  assign n22232 = n7100 & n22231;
  assign n22233 = n7058 & n22232;
  assign n22234 = ~n7057 & n22233;
  assign n22235 = ~n5808 & n22234;
  assign n22236 = ~n6931 & n22235;
  assign n22237 = ~n6056 & n22236;
  assign n22238 = ~n7056 & n22237;
  assign n22239 = n7070 & n22238;
  assign n22240 = n7055 & n22239;
  assign n22241 = n7052 & n22240;
  assign n22242 = ~n22230 & ~n22241;
  assign n22243 = ~n22224 & n22242;
  assign n22244 = n3800 & n19508;
  assign n22245 = n5927 & n22244;
  assign n22246 = n6934 & n22245;
  assign n22247 = ~n6932 & n22246;
  assign n22248 = ~n3940 & n22247;
  assign n22249 = ~n4001 & n22248;
  assign n22250 = ~n5043 & n22249;
  assign n22251 = ~n6931 & n22250;
  assign n22252 = ~n5943 & n22251;
  assign n22253 = ~n6930 & n22252;
  assign n22254 = n6948 & n22253;
  assign n22255 = n6929 & n22254;
  assign n22256 = n6924 & n22255;
  assign n22257 = n7030 & n21161;
  assign n22258 = n7034 & n22257;
  assign n22259 = n6998 & n22258;
  assign n22260 = ~n6997 & n22259;
  assign n22261 = ~n4817 & n22260;
  assign n22262 = ~n4902 & n22261;
  assign n22263 = ~n6931 & n22262;
  assign n22264 = ~n6001 & n22263;
  assign n22265 = ~n6996 & n22264;
  assign n22266 = n7011 & n22265;
  assign n22267 = n6995 & n22266;
  assign n22268 = n6991 & n22267;
  assign n22269 = ~n22256 & ~n22268;
  assign n22270 = pi138 & ~n6432;
  assign n22271 = n7170 & n22270;
  assign n22272 = n7178 & n22271;
  assign n22273 = n6284 & n22272;
  assign n22274 = ~n6784 & n22273;
  assign n22275 = ~n6931 & n22274;
  assign n22276 = ~n6959 & n22275;
  assign n22277 = n7142 & n22276;
  assign n22278 = n7156 & n22277;
  assign n22279 = n7132 & n22278;
  assign n22280 = pi074 & ~n2543;
  assign n22281 = n5772 & n22280;
  assign n22282 = n5776 & n22281;
  assign n22283 = n6875 & n22282;
  assign n22284 = ~n6874 & n22283;
  assign n22285 = ~n3066 & n22284;
  assign n22286 = ~n3983 & n22285;
  assign n22287 = ~n4003 & n22286;
  assign n22288 = ~n4024 & n22287;
  assign n22289 = ~n4999 & n22288;
  assign n22290 = ~n6873 & n22289;
  assign n22291 = ~n5827 & n22290;
  assign n22292 = ~n6872 & n22291;
  assign n22293 = n6890 & n22292;
  assign n22294 = n6871 & n22293;
  assign n22295 = n6866 & n22294;
  assign n22296 = ~n22279 & ~n22295;
  assign n22297 = n22269 & n22296;
  assign n22298 = pi162 & ~n501;
  assign n22299 = n5713 & n22298;
  assign n22300 = n6138 & n22299;
  assign n22301 = n7244 & n22300;
  assign n22302 = ~n1172 & n22301;
  assign n22303 = ~n996 & n22302;
  assign n22304 = ~n2306 & n22303;
  assign n22305 = ~n500 & n22304;
  assign n22306 = n6677 & n22305;
  assign n22307 = n7280 & n22306;
  assign n22308 = n7284 & n22307;
  assign n22309 = ~n7236 & n22308;
  assign n22310 = ~n6137 & n22309;
  assign n22311 = n6193 & n22310;
  assign n22312 = n6134 & n22311;
  assign n22313 = ~n7235 & n22312;
  assign n22314 = n7296 & n22313;
  assign n22315 = n7231 & n22314;
  assign n22316 = ~n6027 & n21131;
  assign n22317 = ~n6931 & n22316;
  assign n22318 = ~n6959 & n22317;
  assign n22319 = n7027 & n22318;
  assign n22320 = n7021 & n22319;
  assign n22321 = ~n6931 & n21182;
  assign n22322 = ~n6114 & n22321;
  assign n22323 = n7054 & n22322;
  assign n22324 = n7093 & n22323;
  assign n22325 = n7087 & n22324;
  assign n22326 = ~n22320 & ~n22325;
  assign n22327 = ~n22315 & n22326;
  assign n22328 = n5835 & n18992;
  assign n22329 = n6843 & n22328;
  assign n22330 = ~n6838 & n22329;
  assign n22331 = ~n2242 & n22330;
  assign n22332 = ~n3095 & n22331;
  assign n22333 = ~n3997 & n22332;
  assign n22334 = ~n4003 & n22333;
  assign n22335 = ~n4837 & n22334;
  assign n22336 = ~n5822 & n22335;
  assign n22337 = ~n6837 & n22336;
  assign n22338 = ~n6820 & n22337;
  assign n22339 = ~n6836 & n22338;
  assign n22340 = n6857 & n22339;
  assign n22341 = n6835 & n22340;
  assign n22342 = n6830 & n22341;
  assign n22343 = ~n5967 & n21109;
  assign n22344 = ~n6931 & n22343;
  assign n22345 = ~n6958 & n22344;
  assign n22346 = n6966 & n22345;
  assign n22347 = ~n5917 & n21112;
  assign n22348 = ~n6911 & n22347;
  assign n22349 = n6916 & n22348;
  assign n22350 = pi154 & ~n501;
  assign n22351 = n7621 & n22350;
  assign n22352 = n7625 & n22351;
  assign n22353 = n7618 & n22352;
  assign n22354 = ~n1172 & n22353;
  assign n22355 = ~n1143 & n22354;
  assign n22356 = ~n996 & n22355;
  assign n22357 = ~n2306 & n22356;
  assign n22358 = ~n500 & n22357;
  assign n22359 = n2316 & n22358;
  assign n22360 = n7608 & n22359;
  assign n22361 = n7757 & n22360;
  assign n22362 = n21848 & n22361;
  assign n22363 = n7597 & n22362;
  assign n22364 = ~n6137 & n22363;
  assign n22365 = n6193 & n22364;
  assign n22366 = n6134 & n22365;
  assign n22367 = ~n22349 & ~n22366;
  assign n22368 = ~n22346 & n22367;
  assign n22369 = ~n22342 & n22368;
  assign n22370 = n22327 & n22369;
  assign n22371 = n22297 & n22370;
  assign po083 = ~n22243 | ~n22371;
  assign n22373 = ~n1026 & n21216;
  assign n22374 = n6787 & n22373;
  assign n22375 = n1239 & n22374;
  assign n22376 = ~n1270 & n22375;
  assign n22377 = n844 & n22376;
  assign n22378 = ~n1372 & n22377;
  assign n22379 = ~n2243 & n22378;
  assign n22380 = ~n6785 & n22379;
  assign n22381 = ~n3104 & n22380;
  assign n22382 = ~n3971 & n22381;
  assign n22383 = ~n4003 & n22382;
  assign n22384 = ~n4872 & n22383;
  assign n22385 = ~n5801 & n22384;
  assign n22386 = ~n6761 & n22385;
  assign n22387 = ~n6760 & n22386;
  assign n22388 = ~n6759 & n22387;
  assign n22389 = n6822 & n22388;
  assign n22390 = n6758 & n22389;
  assign n22391 = n6722 & n22390;
  assign n22392 = pi147 & ~n7193;
  assign n22393 = ~n6754 & n22392;
  assign n22394 = ~n6931 & n22393;
  assign n22395 = n7054 & n22394;
  assign n22396 = n7202 & n22395;
  assign n22397 = n7192 & n22396;
  assign n22398 = n7096 & n21277;
  assign n22399 = n7100 & n22398;
  assign n22400 = n7058 & n22399;
  assign n22401 = ~n7057 & n22400;
  assign n22402 = ~n5808 & n22401;
  assign n22403 = ~n6931 & n22402;
  assign n22404 = ~n6056 & n22403;
  assign n22405 = ~n7056 & n22404;
  assign n22406 = n7070 & n22405;
  assign n22407 = n7055 & n22406;
  assign n22408 = n7052 & n22407;
  assign n22409 = ~n22397 & ~n22408;
  assign n22410 = ~n22391 & n22409;
  assign n22411 = n3800 & n19579;
  assign n22412 = n5927 & n22411;
  assign n22413 = n6934 & n22412;
  assign n22414 = ~n6932 & n22413;
  assign n22415 = ~n3940 & n22414;
  assign n22416 = ~n4001 & n22415;
  assign n22417 = ~n5043 & n22416;
  assign n22418 = ~n6931 & n22417;
  assign n22419 = ~n5943 & n22418;
  assign n22420 = ~n6930 & n22419;
  assign n22421 = n6948 & n22420;
  assign n22422 = n6929 & n22421;
  assign n22423 = n6924 & n22422;
  assign n22424 = n7030 & n21287;
  assign n22425 = n7034 & n22424;
  assign n22426 = n6998 & n22425;
  assign n22427 = ~n6997 & n22426;
  assign n22428 = ~n4817 & n22427;
  assign n22429 = ~n4902 & n22428;
  assign n22430 = ~n6931 & n22429;
  assign n22431 = ~n6001 & n22430;
  assign n22432 = ~n6996 & n22431;
  assign n22433 = n7011 & n22432;
  assign n22434 = n6995 & n22433;
  assign n22435 = n6991 & n22434;
  assign n22436 = ~n22423 & ~n22435;
  assign n22437 = pi139 & ~n6432;
  assign n22438 = n7170 & n22437;
  assign n22439 = n7178 & n22438;
  assign n22440 = n6284 & n22439;
  assign n22441 = ~n6784 & n22440;
  assign n22442 = ~n6931 & n22441;
  assign n22443 = ~n6959 & n22442;
  assign n22444 = n7142 & n22443;
  assign n22445 = n7156 & n22444;
  assign n22446 = n7132 & n22445;
  assign n22447 = pi075 & ~n2543;
  assign n22448 = n5772 & n22447;
  assign n22449 = n5776 & n22448;
  assign n22450 = n6875 & n22449;
  assign n22451 = ~n6874 & n22450;
  assign n22452 = ~n3066 & n22451;
  assign n22453 = ~n3983 & n22452;
  assign n22454 = ~n4003 & n22453;
  assign n22455 = ~n4024 & n22454;
  assign n22456 = ~n4999 & n22455;
  assign n22457 = ~n6873 & n22456;
  assign n22458 = ~n5827 & n22457;
  assign n22459 = ~n6872 & n22458;
  assign n22460 = n6890 & n22459;
  assign n22461 = n6871 & n22460;
  assign n22462 = n6866 & n22461;
  assign n22463 = ~n22446 & ~n22462;
  assign n22464 = n22436 & n22463;
  assign n22465 = pi163 & ~n501;
  assign n22466 = n5713 & n22465;
  assign n22467 = n6138 & n22466;
  assign n22468 = n7244 & n22467;
  assign n22469 = ~n1172 & n22468;
  assign n22470 = ~n996 & n22469;
  assign n22471 = ~n2306 & n22470;
  assign n22472 = ~n500 & n22471;
  assign n22473 = n6677 & n22472;
  assign n22474 = n7280 & n22473;
  assign n22475 = n7284 & n22474;
  assign n22476 = ~n7236 & n22475;
  assign n22477 = ~n6137 & n22476;
  assign n22478 = n6193 & n22477;
  assign n22479 = n6134 & n22478;
  assign n22480 = ~n7235 & n22479;
  assign n22481 = n7296 & n22480;
  assign n22482 = n7231 & n22481;
  assign n22483 = ~n6027 & n21257;
  assign n22484 = ~n6931 & n22483;
  assign n22485 = ~n6959 & n22484;
  assign n22486 = n7027 & n22485;
  assign n22487 = n7021 & n22486;
  assign n22488 = ~n6931 & n21308;
  assign n22489 = ~n6114 & n22488;
  assign n22490 = n7054 & n22489;
  assign n22491 = n7093 & n22490;
  assign n22492 = n7087 & n22491;
  assign n22493 = ~n22487 & ~n22492;
  assign n22494 = ~n22482 & n22493;
  assign n22495 = n5835 & n19051;
  assign n22496 = n6843 & n22495;
  assign n22497 = ~n6838 & n22496;
  assign n22498 = ~n2242 & n22497;
  assign n22499 = ~n3095 & n22498;
  assign n22500 = ~n3997 & n22499;
  assign n22501 = ~n4003 & n22500;
  assign n22502 = ~n4837 & n22501;
  assign n22503 = ~n5822 & n22502;
  assign n22504 = ~n6837 & n22503;
  assign n22505 = ~n6820 & n22504;
  assign n22506 = ~n6836 & n22505;
  assign n22507 = n6857 & n22506;
  assign n22508 = n6835 & n22507;
  assign n22509 = n6830 & n22508;
  assign n22510 = ~n5967 & n21235;
  assign n22511 = ~n6931 & n22510;
  assign n22512 = ~n6958 & n22511;
  assign n22513 = n6966 & n22512;
  assign n22514 = ~n5917 & n21238;
  assign n22515 = ~n6911 & n22514;
  assign n22516 = n6916 & n22515;
  assign n22517 = pi155 & ~n501;
  assign n22518 = n7621 & n22517;
  assign n22519 = n7625 & n22518;
  assign n22520 = n7618 & n22519;
  assign n22521 = ~n1172 & n22520;
  assign n22522 = ~n1143 & n22521;
  assign n22523 = ~n996 & n22522;
  assign n22524 = ~n2306 & n22523;
  assign n22525 = ~n500 & n22524;
  assign n22526 = n2316 & n22525;
  assign n22527 = n7608 & n22526;
  assign n22528 = n7757 & n22527;
  assign n22529 = n21848 & n22528;
  assign n22530 = n7597 & n22529;
  assign n22531 = ~n6137 & n22530;
  assign n22532 = n6193 & n22531;
  assign n22533 = n6134 & n22532;
  assign n22534 = ~n22516 & ~n22533;
  assign n22535 = ~n22513 & n22534;
  assign n22536 = ~n22509 & n22535;
  assign n22537 = n22494 & n22536;
  assign n22538 = n22464 & n22537;
  assign po084 = ~n22410 | ~n22538;
  assign n22540 = ~n1026 & n21342;
  assign n22541 = n6787 & n22540;
  assign n22542 = n1239 & n22541;
  assign n22543 = ~n1270 & n22542;
  assign n22544 = n844 & n22543;
  assign n22545 = ~n1372 & n22544;
  assign n22546 = ~n2243 & n22545;
  assign n22547 = ~n6785 & n22546;
  assign n22548 = ~n3104 & n22547;
  assign n22549 = ~n3971 & n22548;
  assign n22550 = ~n4003 & n22549;
  assign n22551 = ~n4872 & n22550;
  assign n22552 = ~n5801 & n22551;
  assign n22553 = ~n6761 & n22552;
  assign n22554 = ~n6760 & n22553;
  assign n22555 = ~n6759 & n22554;
  assign n22556 = n6822 & n22555;
  assign n22557 = n6758 & n22556;
  assign n22558 = n6722 & n22557;
  assign n22559 = pi148 & ~n7193;
  assign n22560 = ~n6754 & n22559;
  assign n22561 = ~n6931 & n22560;
  assign n22562 = n7054 & n22561;
  assign n22563 = n7202 & n22562;
  assign n22564 = n7192 & n22563;
  assign n22565 = n7096 & n21403;
  assign n22566 = n7100 & n22565;
  assign n22567 = n7058 & n22566;
  assign n22568 = ~n7057 & n22567;
  assign n22569 = ~n5808 & n22568;
  assign n22570 = ~n6931 & n22569;
  assign n22571 = ~n6056 & n22570;
  assign n22572 = ~n7056 & n22571;
  assign n22573 = n7070 & n22572;
  assign n22574 = n7055 & n22573;
  assign n22575 = n7052 & n22574;
  assign n22576 = ~n22564 & ~n22575;
  assign n22577 = ~n22558 & n22576;
  assign n22578 = n3800 & n19650;
  assign n22579 = n5927 & n22578;
  assign n22580 = n6934 & n22579;
  assign n22581 = ~n6932 & n22580;
  assign n22582 = ~n3940 & n22581;
  assign n22583 = ~n4001 & n22582;
  assign n22584 = ~n5043 & n22583;
  assign n22585 = ~n6931 & n22584;
  assign n22586 = ~n5943 & n22585;
  assign n22587 = ~n6930 & n22586;
  assign n22588 = n6948 & n22587;
  assign n22589 = n6929 & n22588;
  assign n22590 = n6924 & n22589;
  assign n22591 = n7030 & n21413;
  assign n22592 = n7034 & n22591;
  assign n22593 = n6998 & n22592;
  assign n22594 = ~n6997 & n22593;
  assign n22595 = ~n4817 & n22594;
  assign n22596 = ~n4902 & n22595;
  assign n22597 = ~n6931 & n22596;
  assign n22598 = ~n6001 & n22597;
  assign n22599 = ~n6996 & n22598;
  assign n22600 = n7011 & n22599;
  assign n22601 = n6995 & n22600;
  assign n22602 = n6991 & n22601;
  assign n22603 = ~n22590 & ~n22602;
  assign n22604 = pi140 & ~n6432;
  assign n22605 = n7170 & n22604;
  assign n22606 = n7178 & n22605;
  assign n22607 = n6284 & n22606;
  assign n22608 = ~n6784 & n22607;
  assign n22609 = ~n6931 & n22608;
  assign n22610 = ~n6959 & n22609;
  assign n22611 = n7142 & n22610;
  assign n22612 = n7156 & n22611;
  assign n22613 = n7132 & n22612;
  assign n22614 = pi076 & ~n2543;
  assign n22615 = n5772 & n22614;
  assign n22616 = n5776 & n22615;
  assign n22617 = n6875 & n22616;
  assign n22618 = ~n6874 & n22617;
  assign n22619 = ~n3066 & n22618;
  assign n22620 = ~n3983 & n22619;
  assign n22621 = ~n4003 & n22620;
  assign n22622 = ~n4024 & n22621;
  assign n22623 = ~n4999 & n22622;
  assign n22624 = ~n6873 & n22623;
  assign n22625 = ~n5827 & n22624;
  assign n22626 = ~n6872 & n22625;
  assign n22627 = n6890 & n22626;
  assign n22628 = n6871 & n22627;
  assign n22629 = n6866 & n22628;
  assign n22630 = ~n22613 & ~n22629;
  assign n22631 = n22603 & n22630;
  assign n22632 = pi164 & ~n501;
  assign n22633 = n5713 & n22632;
  assign n22634 = n6138 & n22633;
  assign n22635 = n7244 & n22634;
  assign n22636 = ~n1172 & n22635;
  assign n22637 = ~n996 & n22636;
  assign n22638 = ~n2306 & n22637;
  assign n22639 = ~n500 & n22638;
  assign n22640 = n6677 & n22639;
  assign n22641 = n7280 & n22640;
  assign n22642 = n7284 & n22641;
  assign n22643 = ~n7236 & n22642;
  assign n22644 = ~n6137 & n22643;
  assign n22645 = n6193 & n22644;
  assign n22646 = n6134 & n22645;
  assign n22647 = ~n7235 & n22646;
  assign n22648 = n7296 & n22647;
  assign n22649 = n7231 & n22648;
  assign n22650 = ~n6027 & n21383;
  assign n22651 = ~n6931 & n22650;
  assign n22652 = ~n6959 & n22651;
  assign n22653 = n7027 & n22652;
  assign n22654 = n7021 & n22653;
  assign n22655 = ~n6931 & n21434;
  assign n22656 = ~n6114 & n22655;
  assign n22657 = n7054 & n22656;
  assign n22658 = n7093 & n22657;
  assign n22659 = n7087 & n22658;
  assign n22660 = ~n22654 & ~n22659;
  assign n22661 = ~n22649 & n22660;
  assign n22662 = n5835 & n19110;
  assign n22663 = n6843 & n22662;
  assign n22664 = ~n6838 & n22663;
  assign n22665 = ~n2242 & n22664;
  assign n22666 = ~n3095 & n22665;
  assign n22667 = ~n3997 & n22666;
  assign n22668 = ~n4003 & n22667;
  assign n22669 = ~n4837 & n22668;
  assign n22670 = ~n5822 & n22669;
  assign n22671 = ~n6837 & n22670;
  assign n22672 = ~n6820 & n22671;
  assign n22673 = ~n6836 & n22672;
  assign n22674 = n6857 & n22673;
  assign n22675 = n6835 & n22674;
  assign n22676 = n6830 & n22675;
  assign n22677 = ~n5967 & n21361;
  assign n22678 = ~n6931 & n22677;
  assign n22679 = ~n6958 & n22678;
  assign n22680 = n6966 & n22679;
  assign n22681 = ~n5917 & n21364;
  assign n22682 = ~n6911 & n22681;
  assign n22683 = n6916 & n22682;
  assign n22684 = pi156 & ~n501;
  assign n22685 = n7621 & n22684;
  assign n22686 = n7625 & n22685;
  assign n22687 = n7618 & n22686;
  assign n22688 = ~n1172 & n22687;
  assign n22689 = ~n1143 & n22688;
  assign n22690 = ~n996 & n22689;
  assign n22691 = ~n2306 & n22690;
  assign n22692 = ~n500 & n22691;
  assign n22693 = n2316 & n22692;
  assign n22694 = n7608 & n22693;
  assign n22695 = n7757 & n22694;
  assign n22696 = n21848 & n22695;
  assign n22697 = n7597 & n22696;
  assign n22698 = ~n6137 & n22697;
  assign n22699 = n6193 & n22698;
  assign n22700 = n6134 & n22699;
  assign n22701 = ~n22683 & ~n22700;
  assign n22702 = ~n22680 & n22701;
  assign n22703 = ~n22676 & n22702;
  assign n22704 = n22661 & n22703;
  assign n22705 = n22631 & n22704;
  assign po085 = ~n22577 | ~n22705;
  assign n22707 = ~n1026 & n21468;
  assign n22708 = n6787 & n22707;
  assign n22709 = n1239 & n22708;
  assign n22710 = ~n1270 & n22709;
  assign n22711 = n844 & n22710;
  assign n22712 = ~n1372 & n22711;
  assign n22713 = ~n2243 & n22712;
  assign n22714 = ~n6785 & n22713;
  assign n22715 = ~n3104 & n22714;
  assign n22716 = ~n3971 & n22715;
  assign n22717 = ~n4003 & n22716;
  assign n22718 = ~n4872 & n22717;
  assign n22719 = ~n5801 & n22718;
  assign n22720 = ~n6761 & n22719;
  assign n22721 = ~n6760 & n22720;
  assign n22722 = ~n6759 & n22721;
  assign n22723 = n6822 & n22722;
  assign n22724 = n6758 & n22723;
  assign n22725 = n6722 & n22724;
  assign n22726 = pi149 & ~n7193;
  assign n22727 = ~n6754 & n22726;
  assign n22728 = ~n6931 & n22727;
  assign n22729 = n7054 & n22728;
  assign n22730 = n7202 & n22729;
  assign n22731 = n7192 & n22730;
  assign n22732 = n7096 & n21529;
  assign n22733 = n7100 & n22732;
  assign n22734 = n7058 & n22733;
  assign n22735 = ~n7057 & n22734;
  assign n22736 = ~n5808 & n22735;
  assign n22737 = ~n6931 & n22736;
  assign n22738 = ~n6056 & n22737;
  assign n22739 = ~n7056 & n22738;
  assign n22740 = n7070 & n22739;
  assign n22741 = n7055 & n22740;
  assign n22742 = n7052 & n22741;
  assign n22743 = ~n22731 & ~n22742;
  assign n22744 = ~n22725 & n22743;
  assign n22745 = n3800 & n19721;
  assign n22746 = n5927 & n22745;
  assign n22747 = n6934 & n22746;
  assign n22748 = ~n6932 & n22747;
  assign n22749 = ~n3940 & n22748;
  assign n22750 = ~n4001 & n22749;
  assign n22751 = ~n5043 & n22750;
  assign n22752 = ~n6931 & n22751;
  assign n22753 = ~n5943 & n22752;
  assign n22754 = ~n6930 & n22753;
  assign n22755 = n6948 & n22754;
  assign n22756 = n6929 & n22755;
  assign n22757 = n6924 & n22756;
  assign n22758 = n7030 & n21539;
  assign n22759 = n7034 & n22758;
  assign n22760 = n6998 & n22759;
  assign n22761 = ~n6997 & n22760;
  assign n22762 = ~n4817 & n22761;
  assign n22763 = ~n4902 & n22762;
  assign n22764 = ~n6931 & n22763;
  assign n22765 = ~n6001 & n22764;
  assign n22766 = ~n6996 & n22765;
  assign n22767 = n7011 & n22766;
  assign n22768 = n6995 & n22767;
  assign n22769 = n6991 & n22768;
  assign n22770 = ~n22757 & ~n22769;
  assign n22771 = pi141 & ~n6432;
  assign n22772 = n7170 & n22771;
  assign n22773 = n7178 & n22772;
  assign n22774 = n6284 & n22773;
  assign n22775 = ~n6784 & n22774;
  assign n22776 = ~n6931 & n22775;
  assign n22777 = ~n6959 & n22776;
  assign n22778 = n7142 & n22777;
  assign n22779 = n7156 & n22778;
  assign n22780 = n7132 & n22779;
  assign n22781 = pi077 & ~n2543;
  assign n22782 = n5772 & n22781;
  assign n22783 = n5776 & n22782;
  assign n22784 = n6875 & n22783;
  assign n22785 = ~n6874 & n22784;
  assign n22786 = ~n3066 & n22785;
  assign n22787 = ~n3983 & n22786;
  assign n22788 = ~n4003 & n22787;
  assign n22789 = ~n4024 & n22788;
  assign n22790 = ~n4999 & n22789;
  assign n22791 = ~n6873 & n22790;
  assign n22792 = ~n5827 & n22791;
  assign n22793 = ~n6872 & n22792;
  assign n22794 = n6890 & n22793;
  assign n22795 = n6871 & n22794;
  assign n22796 = n6866 & n22795;
  assign n22797 = ~n22780 & ~n22796;
  assign n22798 = n22770 & n22797;
  assign n22799 = pi165 & ~n501;
  assign n22800 = n5713 & n22799;
  assign n22801 = n6138 & n22800;
  assign n22802 = n7244 & n22801;
  assign n22803 = ~n1172 & n22802;
  assign n22804 = ~n996 & n22803;
  assign n22805 = ~n2306 & n22804;
  assign n22806 = ~n500 & n22805;
  assign n22807 = n6677 & n22806;
  assign n22808 = n7280 & n22807;
  assign n22809 = n7284 & n22808;
  assign n22810 = ~n7236 & n22809;
  assign n22811 = ~n6137 & n22810;
  assign n22812 = n6193 & n22811;
  assign n22813 = n6134 & n22812;
  assign n22814 = ~n7235 & n22813;
  assign n22815 = n7296 & n22814;
  assign n22816 = n7231 & n22815;
  assign n22817 = ~n6027 & n21509;
  assign n22818 = ~n6931 & n22817;
  assign n22819 = ~n6959 & n22818;
  assign n22820 = n7027 & n22819;
  assign n22821 = n7021 & n22820;
  assign n22822 = ~n6931 & n21560;
  assign n22823 = ~n6114 & n22822;
  assign n22824 = n7054 & n22823;
  assign n22825 = n7093 & n22824;
  assign n22826 = n7087 & n22825;
  assign n22827 = ~n22821 & ~n22826;
  assign n22828 = ~n22816 & n22827;
  assign n22829 = n5835 & n19169;
  assign n22830 = n6843 & n22829;
  assign n22831 = ~n6838 & n22830;
  assign n22832 = ~n2242 & n22831;
  assign n22833 = ~n3095 & n22832;
  assign n22834 = ~n3997 & n22833;
  assign n22835 = ~n4003 & n22834;
  assign n22836 = ~n4837 & n22835;
  assign n22837 = ~n5822 & n22836;
  assign n22838 = ~n6837 & n22837;
  assign n22839 = ~n6820 & n22838;
  assign n22840 = ~n6836 & n22839;
  assign n22841 = n6857 & n22840;
  assign n22842 = n6835 & n22841;
  assign n22843 = n6830 & n22842;
  assign n22844 = ~n5967 & n21487;
  assign n22845 = ~n6931 & n22844;
  assign n22846 = ~n6958 & n22845;
  assign n22847 = n6966 & n22846;
  assign n22848 = ~n5917 & n21490;
  assign n22849 = ~n6911 & n22848;
  assign n22850 = n6916 & n22849;
  assign n22851 = pi157 & ~n501;
  assign n22852 = n7621 & n22851;
  assign n22853 = n7625 & n22852;
  assign n22854 = n7618 & n22853;
  assign n22855 = ~n1172 & n22854;
  assign n22856 = ~n1143 & n22855;
  assign n22857 = ~n996 & n22856;
  assign n22858 = ~n2306 & n22857;
  assign n22859 = ~n500 & n22858;
  assign n22860 = n2316 & n22859;
  assign n22861 = n7608 & n22860;
  assign n22862 = n7757 & n22861;
  assign n22863 = n21848 & n22862;
  assign n22864 = n7597 & n22863;
  assign n22865 = ~n6137 & n22864;
  assign n22866 = n6193 & n22865;
  assign n22867 = n6134 & n22866;
  assign n22868 = ~n22850 & ~n22867;
  assign n22869 = ~n22847 & n22868;
  assign n22870 = ~n22843 & n22869;
  assign n22871 = n22828 & n22870;
  assign n22872 = n22798 & n22871;
  assign po086 = ~n22744 | ~n22872;
  assign n22874 = ~n1026 & n21594;
  assign n22875 = n6787 & n22874;
  assign n22876 = n1239 & n22875;
  assign n22877 = ~n1270 & n22876;
  assign n22878 = n844 & n22877;
  assign n22879 = ~n1372 & n22878;
  assign n22880 = ~n2243 & n22879;
  assign n22881 = ~n6785 & n22880;
  assign n22882 = ~n3104 & n22881;
  assign n22883 = ~n3971 & n22882;
  assign n22884 = ~n4003 & n22883;
  assign n22885 = ~n4872 & n22884;
  assign n22886 = ~n5801 & n22885;
  assign n22887 = ~n6761 & n22886;
  assign n22888 = ~n6760 & n22887;
  assign n22889 = ~n6759 & n22888;
  assign n22890 = n6822 & n22889;
  assign n22891 = n6758 & n22890;
  assign n22892 = n6722 & n22891;
  assign n22893 = pi150 & ~n7193;
  assign n22894 = ~n6754 & n22893;
  assign n22895 = ~n6931 & n22894;
  assign n22896 = n7054 & n22895;
  assign n22897 = n7202 & n22896;
  assign n22898 = n7192 & n22897;
  assign n22899 = n7096 & n21655;
  assign n22900 = n7100 & n22899;
  assign n22901 = n7058 & n22900;
  assign n22902 = ~n7057 & n22901;
  assign n22903 = ~n5808 & n22902;
  assign n22904 = ~n6931 & n22903;
  assign n22905 = ~n6056 & n22904;
  assign n22906 = ~n7056 & n22905;
  assign n22907 = n7070 & n22906;
  assign n22908 = n7055 & n22907;
  assign n22909 = n7052 & n22908;
  assign n22910 = ~n22898 & ~n22909;
  assign n22911 = ~n22892 & n22910;
  assign n22912 = n3800 & n19792;
  assign n22913 = n5927 & n22912;
  assign n22914 = n6934 & n22913;
  assign n22915 = ~n6932 & n22914;
  assign n22916 = ~n3940 & n22915;
  assign n22917 = ~n4001 & n22916;
  assign n22918 = ~n5043 & n22917;
  assign n22919 = ~n6931 & n22918;
  assign n22920 = ~n5943 & n22919;
  assign n22921 = ~n6930 & n22920;
  assign n22922 = n6948 & n22921;
  assign n22923 = n6929 & n22922;
  assign n22924 = n6924 & n22923;
  assign n22925 = n7030 & n21665;
  assign n22926 = n7034 & n22925;
  assign n22927 = n6998 & n22926;
  assign n22928 = ~n6997 & n22927;
  assign n22929 = ~n4817 & n22928;
  assign n22930 = ~n4902 & n22929;
  assign n22931 = ~n6931 & n22930;
  assign n22932 = ~n6001 & n22931;
  assign n22933 = ~n6996 & n22932;
  assign n22934 = n7011 & n22933;
  assign n22935 = n6995 & n22934;
  assign n22936 = n6991 & n22935;
  assign n22937 = ~n22924 & ~n22936;
  assign n22938 = pi142 & ~n6432;
  assign n22939 = n7170 & n22938;
  assign n22940 = n7178 & n22939;
  assign n22941 = n6284 & n22940;
  assign n22942 = ~n6784 & n22941;
  assign n22943 = ~n6931 & n22942;
  assign n22944 = ~n6959 & n22943;
  assign n22945 = n7142 & n22944;
  assign n22946 = n7156 & n22945;
  assign n22947 = n7132 & n22946;
  assign n22948 = pi078 & ~n2543;
  assign n22949 = n5772 & n22948;
  assign n22950 = n5776 & n22949;
  assign n22951 = n6875 & n22950;
  assign n22952 = ~n6874 & n22951;
  assign n22953 = ~n3066 & n22952;
  assign n22954 = ~n3983 & n22953;
  assign n22955 = ~n4003 & n22954;
  assign n22956 = ~n4024 & n22955;
  assign n22957 = ~n4999 & n22956;
  assign n22958 = ~n6873 & n22957;
  assign n22959 = ~n5827 & n22958;
  assign n22960 = ~n6872 & n22959;
  assign n22961 = n6890 & n22960;
  assign n22962 = n6871 & n22961;
  assign n22963 = n6866 & n22962;
  assign n22964 = ~n22947 & ~n22963;
  assign n22965 = n22937 & n22964;
  assign n22966 = pi166 & ~n501;
  assign n22967 = n5713 & n22966;
  assign n22968 = n6138 & n22967;
  assign n22969 = n7244 & n22968;
  assign n22970 = ~n1172 & n22969;
  assign n22971 = ~n996 & n22970;
  assign n22972 = ~n2306 & n22971;
  assign n22973 = ~n500 & n22972;
  assign n22974 = n6677 & n22973;
  assign n22975 = n7280 & n22974;
  assign n22976 = n7284 & n22975;
  assign n22977 = ~n7236 & n22976;
  assign n22978 = ~n6137 & n22977;
  assign n22979 = n6193 & n22978;
  assign n22980 = n6134 & n22979;
  assign n22981 = ~n7235 & n22980;
  assign n22982 = n7296 & n22981;
  assign n22983 = n7231 & n22982;
  assign n22984 = ~n6027 & n21635;
  assign n22985 = ~n6931 & n22984;
  assign n22986 = ~n6959 & n22985;
  assign n22987 = n7027 & n22986;
  assign n22988 = n7021 & n22987;
  assign n22989 = ~n6931 & n21686;
  assign n22990 = ~n6114 & n22989;
  assign n22991 = n7054 & n22990;
  assign n22992 = n7093 & n22991;
  assign n22993 = n7087 & n22992;
  assign n22994 = ~n22988 & ~n22993;
  assign n22995 = ~n22983 & n22994;
  assign n22996 = n5835 & n19228;
  assign n22997 = n6843 & n22996;
  assign n22998 = ~n6838 & n22997;
  assign n22999 = ~n2242 & n22998;
  assign n23000 = ~n3095 & n22999;
  assign n23001 = ~n3997 & n23000;
  assign n23002 = ~n4003 & n23001;
  assign n23003 = ~n4837 & n23002;
  assign n23004 = ~n5822 & n23003;
  assign n23005 = ~n6837 & n23004;
  assign n23006 = ~n6820 & n23005;
  assign n23007 = ~n6836 & n23006;
  assign n23008 = n6857 & n23007;
  assign n23009 = n6835 & n23008;
  assign n23010 = n6830 & n23009;
  assign n23011 = ~n5967 & n21613;
  assign n23012 = ~n6931 & n23011;
  assign n23013 = ~n6958 & n23012;
  assign n23014 = n6966 & n23013;
  assign n23015 = ~n5917 & n21616;
  assign n23016 = ~n6911 & n23015;
  assign n23017 = n6916 & n23016;
  assign n23018 = pi158 & ~n501;
  assign n23019 = n7621 & n23018;
  assign n23020 = n7625 & n23019;
  assign n23021 = n7618 & n23020;
  assign n23022 = ~n1172 & n23021;
  assign n23023 = ~n1143 & n23022;
  assign n23024 = ~n996 & n23023;
  assign n23025 = ~n2306 & n23024;
  assign n23026 = ~n500 & n23025;
  assign n23027 = n2316 & n23026;
  assign n23028 = n7608 & n23027;
  assign n23029 = n7757 & n23028;
  assign n23030 = n21848 & n23029;
  assign n23031 = n7597 & n23030;
  assign n23032 = ~n6137 & n23031;
  assign n23033 = n6193 & n23032;
  assign n23034 = n6134 & n23033;
  assign n23035 = ~n23017 & ~n23034;
  assign n23036 = ~n23014 & n23035;
  assign n23037 = ~n23010 & n23036;
  assign n23038 = n22995 & n23037;
  assign n23039 = n22965 & n23038;
  assign po087 = ~n22911 | ~n23039;
  assign n23041 = ~n6967 & n21792;
  assign n23042 = ~n8017 & n23041;
  assign n23043 = ~n8044 & n23042;
  assign n23044 = n8052 & n23043;
  assign n23045 = pi175 & ~n501;
  assign n23046 = n5714 & n23045;
  assign n23047 = n5719 & n23046;
  assign n23048 = n8912 & n23047;
  assign n23049 = ~n1172 & n23048;
  assign n23050 = ~n996 & n23049;
  assign n23051 = ~n2306 & n23050;
  assign n23052 = ~n500 & n23051;
  assign n23053 = n6677 & n23052;
  assign n23054 = n8880 & n23053;
  assign n23055 = n7284 & n23054;
  assign n23056 = ~n7236 & n23055;
  assign n23057 = ~n6137 & n23056;
  assign n23058 = n6193 & n23057;
  assign n23059 = n6134 & n23058;
  assign n23060 = ~n8867 & n23059;
  assign n23061 = ~n7235 & n23060;
  assign n23062 = n7296 & n23061;
  assign n23063 = n7231 & n23062;
  assign n23064 = ~n8866 & n23063;
  assign n23065 = n8898 & n23064;
  assign n23066 = n8863 & n23065;
  assign n23067 = ~n7029 & n21796;
  assign n23068 = ~n8017 & n23067;
  assign n23069 = ~n8045 & n23068;
  assign n23070 = n8143 & n23069;
  assign n23071 = n8137 & n23070;
  assign n23072 = ~n23066 & ~n23071;
  assign n23073 = ~n23044 & n23072;
  assign n23074 = n3740 & n20682;
  assign n23075 = n3951 & n23074;
  assign n23076 = n3680 & n4100;
  assign n23077 = ~n3464 & n23076;
  assign n23078 = ~n3165 & n23077;
  assign n23079 = n23075 & n23078;
  assign n23080 = ~n3940 & n23079;
  assign n23081 = ~n4001 & n23080;
  assign n23082 = ~n5043 & n23081;
  assign n23083 = ~n5943 & n23082;
  assign n23084 = ~n8018 & n23083;
  assign n23085 = ~n8017 & n23084;
  assign n23086 = ~n6951 & n23085;
  assign n23087 = ~n8016 & n23086;
  assign n23088 = n8034 & n23087;
  assign n23089 = n8015 & n23088;
  assign n23090 = n8008 & n23089;
  assign n23091 = ~n6114 & n20804;
  assign n23092 = ~n7095 & n23091;
  assign n23093 = ~n8017 & n23092;
  assign n23094 = n8155 & n23093;
  assign n23095 = n8216 & n23094;
  assign n23096 = n8210 & n23095;
  assign n23097 = ~n6917 & n21841;
  assign n23098 = ~n7993 & n23097;
  assign n23099 = n7998 & n23098;
  assign n23100 = pi167 & ~n501;
  assign n23101 = n8692 & n23100;
  assign n23102 = n8941 & n23101;
  assign n23103 = n8946 & n23102;
  assign n23104 = n8940 & n23103;
  assign n23105 = ~n1172 & n23104;
  assign n23106 = ~n1025 & n23105;
  assign n23107 = ~n996 & n23106;
  assign n23108 = n8701 & n23107;
  assign n23109 = n3821 & n23108;
  assign n23110 = n8681 & n23109;
  assign n23111 = n8824 & n23110;
  assign n23112 = n8679 & n23111;
  assign n23113 = n8666 & n23112;
  assign n23114 = ~n7236 & n23113;
  assign n23115 = ~n6137 & n23114;
  assign n23116 = n6193 & n23115;
  assign n23117 = n6134 & n23116;
  assign n23118 = ~n7235 & n23117;
  assign n23119 = n7296 & n23118;
  assign n23120 = n7231 & n23119;
  assign n23121 = ~n23099 & ~n23120;
  assign n23122 = ~n23096 & n23121;
  assign n23123 = ~n23090 & n23122;
  assign n23124 = n8264 & n21696;
  assign n23125 = ~n6784 & n23124;
  assign n23126 = ~n8232 & n23125;
  assign n23127 = ~n8017 & n23126;
  assign n23128 = ~n7158 & n23127;
  assign n23129 = ~n8231 & n23128;
  assign n23130 = n8247 & n23129;
  assign n23131 = n8230 & n23130;
  assign n23132 = n8227 & n23131;
  assign n23133 = pi151 & ~n7659;
  assign n23134 = ~n7660 & n23133;
  assign n23135 = ~n7658 & n23134;
  assign n23136 = ~n7692 & n23135;
  assign n23137 = n7752 & n23136;
  assign n23138 = n7536 & n23137;
  assign n23139 = n8338 & n23138;
  assign n23140 = ~n7869 & n23139;
  assign n23141 = ~n8017 & n23140;
  assign n23142 = ~n8045 & n23141;
  assign n23143 = ~n8335 & n23142;
  assign n23144 = n8331 & n23143;
  assign n23145 = n8328 & n23144;
  assign n23146 = n8306 & n23145;
  assign n23147 = ~n23132 & ~n23146;
  assign n23148 = n23123 & n23147;
  assign n23149 = n23073 & n23148;
  assign n23150 = n8121 & n21731;
  assign n23151 = ~n4817 & n23150;
  assign n23152 = ~n4902 & n23151;
  assign n23153 = ~n6001 & n23152;
  assign n23154 = ~n8094 & n23153;
  assign n23155 = ~n8017 & n23154;
  assign n23156 = ~n7014 & n23155;
  assign n23157 = ~n8093 & n23156;
  assign n23158 = n8111 & n23157;
  assign n23159 = n8092 & n23158;
  assign n23160 = n8086 & n23159;
  assign n23161 = pi143 & ~n6754;
  assign n23162 = ~n8017 & n23161;
  assign n23163 = ~n7204 & n23162;
  assign n23164 = ~n8282 & n23163;
  assign n23165 = n8288 & n23164;
  assign n23166 = n8281 & n23165;
  assign n23167 = n8280 & n23166;
  assign n23168 = n3846 & n21711;
  assign n23169 = n3854 & n23168;
  assign n23170 = n3849 & n7974;
  assign n23171 = ~n3024 & n23170;
  assign n23172 = ~n2934 & n23171;
  assign n23173 = n23169 & n23172;
  assign n23174 = ~n3066 & n23173;
  assign n23175 = ~n3983 & n23174;
  assign n23176 = ~n4003 & n23175;
  assign n23177 = ~n4024 & n23176;
  assign n23178 = ~n4999 & n23177;
  assign n23179 = ~n5827 & n23178;
  assign n23180 = ~n7870 & n23179;
  assign n23181 = ~n7842 & n23180;
  assign n23182 = ~n6893 & n23181;
  assign n23183 = ~n7841 & n23182;
  assign n23184 = n7887 & n23183;
  assign n23185 = n7840 & n23184;
  assign n23186 = n7810 & n23185;
  assign n23187 = ~n23167 & ~n23186;
  assign n23188 = ~n23160 & n23187;
  assign n23189 = ~n5524 & n20770;
  assign n23190 = ~n5522 & n23189;
  assign n23191 = ~n5598 & n23190;
  assign n23192 = n6068 & n23191;
  assign n23193 = n6066 & n23192;
  assign n23194 = ~n5469 & n6075;
  assign n23195 = ~n5170 & n23194;
  assign n23196 = n23193 & n23195;
  assign n23197 = ~n5808 & n23196;
  assign n23198 = ~n6056 & n23197;
  assign n23199 = ~n8161 & n23198;
  assign n23200 = ~n8017 & n23199;
  assign n23201 = ~n7073 & n23200;
  assign n23202 = ~n8160 & n23201;
  assign n23203 = n8176 & n23202;
  assign n23204 = n8159 & n23203;
  assign n23205 = n8154 & n23204;
  assign n23206 = pi039 & ~n1115;
  assign n23207 = ~n1026 & n23206;
  assign n23208 = ~n1086 & n23207;
  assign n23209 = n1239 & n23208;
  assign n23210 = ~n1270 & n23209;
  assign n23211 = n844 & n23210;
  assign n23212 = ~n1372 & n23211;
  assign n23213 = ~n2243 & n23212;
  assign n23214 = ~n3104 & n23213;
  assign n23215 = ~n3971 & n23214;
  assign n23216 = ~n4003 & n23215;
  assign n23217 = ~n4872 & n23216;
  assign n23218 = ~n5801 & n23217;
  assign n23219 = ~n6739 & n23218;
  assign n23220 = ~n7945 & n23219;
  assign n23221 = ~n7944 & n23220;
  assign n23222 = ~n7807 & n23221;
  assign n23223 = ~n7943 & n23222;
  assign n23224 = n7966 & n23223;
  assign n23225 = n7942 & n23224;
  assign n23226 = n7935 & n23225;
  assign n23227 = ~n23205 & ~n23226;
  assign n23228 = pi159 & ~n8391;
  assign n23229 = ~po161 & n23228;
  assign n23230 = ~n8017 & n23229;
  assign n23231 = ~n8314 & n23230;
  assign n23232 = n8281 & n23231;
  assign n23233 = n8390 & n23232;
  assign n23234 = n8383 & n23233;
  assign n23235 = ~n1958 & n18802;
  assign n23236 = n7910 & n23235;
  assign n23237 = ~n2242 & n23236;
  assign n23238 = ~n3095 & n23237;
  assign n23239 = ~n3997 & n23238;
  assign n23240 = ~n4003 & n23239;
  assign n23241 = ~n4837 & n23240;
  assign n23242 = ~n5822 & n23241;
  assign n23243 = ~n6820 & n23242;
  assign n23244 = ~n7907 & n23243;
  assign n23245 = ~n7906 & n23244;
  assign n23246 = ~n7785 & n23245;
  assign n23247 = ~n7905 & n23246;
  assign n23248 = n7925 & n23247;
  assign n23249 = n7904 & n23248;
  assign n23250 = n7897 & n23249;
  assign n23251 = ~n23234 & ~n23250;
  assign n23252 = n23227 & n23251;
  assign n23253 = n23188 & n23252;
  assign po088 = ~n23149 | ~n23253;
  assign n23255 = ~n6967 & n21970;
  assign n23256 = ~n8017 & n23255;
  assign n23257 = ~n8044 & n23256;
  assign n23258 = n8052 & n23257;
  assign n23259 = ~n6114 & n20919;
  assign n23260 = ~n7095 & n23259;
  assign n23261 = ~n8017 & n23260;
  assign n23262 = n8155 & n23261;
  assign n23263 = n8216 & n23262;
  assign n23264 = n8210 & n23263;
  assign n23265 = pi176 & ~n501;
  assign n23266 = n5714 & n23265;
  assign n23267 = n5719 & n23266;
  assign n23268 = n8912 & n23267;
  assign n23269 = ~n1172 & n23268;
  assign n23270 = ~n996 & n23269;
  assign n23271 = ~n2306 & n23270;
  assign n23272 = ~n500 & n23271;
  assign n23273 = n6677 & n23272;
  assign n23274 = n8880 & n23273;
  assign n23275 = n7284 & n23274;
  assign n23276 = ~n7236 & n23275;
  assign n23277 = ~n6137 & n23276;
  assign n23278 = n6193 & n23277;
  assign n23279 = n6134 & n23278;
  assign n23280 = ~n8867 & n23279;
  assign n23281 = ~n7235 & n23280;
  assign n23282 = n7296 & n23281;
  assign n23283 = n7231 & n23282;
  assign n23284 = ~n8866 & n23283;
  assign n23285 = n8898 & n23284;
  assign n23286 = n8863 & n23285;
  assign n23287 = ~n23264 & ~n23286;
  assign n23288 = ~n23258 & n23287;
  assign n23289 = n8193 & n21872;
  assign n23290 = ~n5808 & n23289;
  assign n23291 = ~n6056 & n23290;
  assign n23292 = ~n8161 & n23291;
  assign n23293 = ~n8017 & n23292;
  assign n23294 = ~n7073 & n23293;
  assign n23295 = ~n8160 & n23294;
  assign n23296 = n8176 & n23295;
  assign n23297 = n8159 & n23296;
  assign n23298 = n8154 & n23297;
  assign n23299 = ~n7029 & n21965;
  assign n23300 = ~n8017 & n23299;
  assign n23301 = ~n8045 & n23300;
  assign n23302 = n8143 & n23301;
  assign n23303 = n8137 & n23302;
  assign n23304 = ~n6917 & n22013;
  assign n23305 = ~n7993 & n23304;
  assign n23306 = n7998 & n23305;
  assign n23307 = pi168 & ~n501;
  assign n23308 = n8692 & n23307;
  assign n23309 = n8941 & n23308;
  assign n23310 = n8946 & n23309;
  assign n23311 = n8940 & n23310;
  assign n23312 = ~n1172 & n23311;
  assign n23313 = ~n1025 & n23312;
  assign n23314 = ~n996 & n23313;
  assign n23315 = n8701 & n23314;
  assign n23316 = n3821 & n23315;
  assign n23317 = n8681 & n23316;
  assign n23318 = n8824 & n23317;
  assign n23319 = n8679 & n23318;
  assign n23320 = n8666 & n23319;
  assign n23321 = ~n7236 & n23320;
  assign n23322 = ~n6137 & n23321;
  assign n23323 = n6193 & n23322;
  assign n23324 = n6134 & n23323;
  assign n23325 = ~n7235 & n23324;
  assign n23326 = n7296 & n23325;
  assign n23327 = n7231 & n23326;
  assign n23328 = ~n23306 & ~n23327;
  assign n23329 = ~n23303 & n23328;
  assign n23330 = ~n23298 & n23329;
  assign n23331 = n8264 & n21949;
  assign n23332 = ~n6784 & n23331;
  assign n23333 = ~n8232 & n23332;
  assign n23334 = ~n8017 & n23333;
  assign n23335 = ~n7158 & n23334;
  assign n23336 = ~n8231 & n23335;
  assign n23337 = n8247 & n23336;
  assign n23338 = n8230 & n23337;
  assign n23339 = n8227 & n23338;
  assign n23340 = n8059 & n21922;
  assign n23341 = ~n3940 & n23340;
  assign n23342 = ~n4001 & n23341;
  assign n23343 = ~n5043 & n23342;
  assign n23344 = ~n5943 & n23343;
  assign n23345 = ~n8018 & n23344;
  assign n23346 = ~n8017 & n23345;
  assign n23347 = ~n6951 & n23346;
  assign n23348 = ~n8016 & n23347;
  assign n23349 = n8034 & n23348;
  assign n23350 = n8015 & n23349;
  assign n23351 = n8008 & n23350;
  assign n23352 = ~n23339 & ~n23351;
  assign n23353 = n23330 & n23352;
  assign n23354 = n23288 & n23353;
  assign n23355 = n8121 & n21936;
  assign n23356 = ~n4817 & n23355;
  assign n23357 = ~n4902 & n23356;
  assign n23358 = ~n6001 & n23357;
  assign n23359 = ~n8094 & n23358;
  assign n23360 = ~n8017 & n23359;
  assign n23361 = ~n7014 & n23360;
  assign n23362 = ~n8093 & n23361;
  assign n23363 = n8111 & n23362;
  assign n23364 = n8092 & n23363;
  assign n23365 = n8086 & n23364;
  assign n23366 = pi040 & ~n1115;
  assign n23367 = ~n1026 & n23366;
  assign n23368 = ~n1086 & n23367;
  assign n23369 = n1239 & n23368;
  assign n23370 = ~n1270 & n23369;
  assign n23371 = n844 & n23370;
  assign n23372 = ~n1372 & n23371;
  assign n23373 = ~n2243 & n23372;
  assign n23374 = ~n3104 & n23373;
  assign n23375 = ~n3971 & n23374;
  assign n23376 = ~n4003 & n23375;
  assign n23377 = ~n4872 & n23376;
  assign n23378 = ~n5801 & n23377;
  assign n23379 = ~n6739 & n23378;
  assign n23380 = ~n7945 & n23379;
  assign n23381 = ~n7944 & n23380;
  assign n23382 = ~n7807 & n23381;
  assign n23383 = ~n7943 & n23382;
  assign n23384 = n7966 & n23383;
  assign n23385 = n7942 & n23384;
  assign n23386 = n7935 & n23385;
  assign n23387 = n7978 & n21884;
  assign n23388 = ~n3066 & n23387;
  assign n23389 = ~n3983 & n23388;
  assign n23390 = ~n4003 & n23389;
  assign n23391 = ~n4024 & n23390;
  assign n23392 = ~n4999 & n23391;
  assign n23393 = ~n5827 & n23392;
  assign n23394 = ~n7870 & n23393;
  assign n23395 = ~n7842 & n23394;
  assign n23396 = ~n6893 & n23395;
  assign n23397 = ~n7841 & n23396;
  assign n23398 = n7887 & n23397;
  assign n23399 = n7840 & n23398;
  assign n23400 = n7810 & n23399;
  assign n23401 = ~n23386 & ~n23400;
  assign n23402 = ~n23365 & n23401;
  assign n23403 = pi152 & ~n7663;
  assign n23404 = n8360 & n23403;
  assign n23405 = n8368 & n23404;
  assign n23406 = ~n7869 & n23405;
  assign n23407 = ~n8017 & n23406;
  assign n23408 = ~n8045 & n23407;
  assign n23409 = ~n8335 & n23408;
  assign n23410 = n8331 & n23409;
  assign n23411 = n8328 & n23410;
  assign n23412 = n8306 & n23411;
  assign n23413 = pi144 & ~n6754;
  assign n23414 = ~n8017 & n23413;
  assign n23415 = ~n7204 & n23414;
  assign n23416 = ~n8282 & n23415;
  assign n23417 = n8288 & n23416;
  assign n23418 = n8281 & n23417;
  assign n23419 = n8280 & n23418;
  assign n23420 = ~n23412 & ~n23419;
  assign n23421 = pi160 & ~n8391;
  assign n23422 = ~po161 & n23421;
  assign n23423 = ~n8017 & n23422;
  assign n23424 = ~n8314 & n23423;
  assign n23425 = n8281 & n23424;
  assign n23426 = n8390 & n23425;
  assign n23427 = n8383 & n23426;
  assign n23428 = ~n1958 & n18861;
  assign n23429 = n7910 & n23428;
  assign n23430 = ~n2242 & n23429;
  assign n23431 = ~n3095 & n23430;
  assign n23432 = ~n3997 & n23431;
  assign n23433 = ~n4003 & n23432;
  assign n23434 = ~n4837 & n23433;
  assign n23435 = ~n5822 & n23434;
  assign n23436 = ~n6820 & n23435;
  assign n23437 = ~n7907 & n23436;
  assign n23438 = ~n7906 & n23437;
  assign n23439 = ~n7785 & n23438;
  assign n23440 = ~n7905 & n23439;
  assign n23441 = n7925 & n23440;
  assign n23442 = n7904 & n23441;
  assign n23443 = n7897 & n23442;
  assign n23444 = ~n23427 & ~n23443;
  assign n23445 = n23420 & n23444;
  assign n23446 = n23402 & n23445;
  assign po089 = ~n23354 | ~n23446;
  assign n23448 = pi177 & ~n501;
  assign n23449 = n5714 & n23448;
  assign n23450 = n5719 & n23449;
  assign n23451 = n8912 & n23450;
  assign n23452 = ~n1172 & n23451;
  assign n23453 = ~n996 & n23452;
  assign n23454 = ~n2306 & n23453;
  assign n23455 = ~n500 & n23454;
  assign n23456 = n6677 & n23455;
  assign n23457 = n8880 & n23456;
  assign n23458 = n7284 & n23457;
  assign n23459 = ~n7236 & n23458;
  assign n23460 = ~n6137 & n23459;
  assign n23461 = n6193 & n23460;
  assign n23462 = n6134 & n23461;
  assign n23463 = ~n8867 & n23462;
  assign n23464 = ~n7235 & n23463;
  assign n23465 = n7296 & n23464;
  assign n23466 = n7231 & n23465;
  assign n23467 = ~n8866 & n23466;
  assign n23468 = n8898 & n23467;
  assign n23469 = n8863 & n23468;
  assign n23470 = ~n7029 & n22151;
  assign n23471 = ~n8017 & n23470;
  assign n23472 = ~n8045 & n23471;
  assign n23473 = n8143 & n23472;
  assign n23474 = n8137 & n23473;
  assign n23475 = ~n6114 & n21056;
  assign n23476 = ~n7095 & n23475;
  assign n23477 = ~n8017 & n23476;
  assign n23478 = n8155 & n23477;
  assign n23479 = n8216 & n23478;
  assign n23480 = n8210 & n23479;
  assign n23481 = ~n23474 & ~n23480;
  assign n23482 = ~n23469 & n23481;
  assign n23483 = n8059 & n22163;
  assign n23484 = ~n3940 & n23483;
  assign n23485 = ~n4001 & n23484;
  assign n23486 = ~n5043 & n23485;
  assign n23487 = ~n5943 & n23486;
  assign n23488 = ~n8018 & n23487;
  assign n23489 = ~n8017 & n23488;
  assign n23490 = ~n6951 & n23489;
  assign n23491 = ~n8016 & n23490;
  assign n23492 = n8034 & n23491;
  assign n23493 = n8015 & n23492;
  assign n23494 = n8008 & n23493;
  assign n23495 = ~n6967 & n22176;
  assign n23496 = ~n8017 & n23495;
  assign n23497 = ~n8044 & n23496;
  assign n23498 = n8052 & n23497;
  assign n23499 = ~n6917 & n22180;
  assign n23500 = ~n7993 & n23499;
  assign n23501 = n7998 & n23500;
  assign n23502 = pi169 & ~n501;
  assign n23503 = n8692 & n23502;
  assign n23504 = n8941 & n23503;
  assign n23505 = n8946 & n23504;
  assign n23506 = n8940 & n23505;
  assign n23507 = ~n1172 & n23506;
  assign n23508 = ~n1025 & n23507;
  assign n23509 = ~n996 & n23508;
  assign n23510 = n8701 & n23509;
  assign n23511 = n3821 & n23510;
  assign n23512 = n8681 & n23511;
  assign n23513 = n8824 & n23512;
  assign n23514 = n8679 & n23513;
  assign n23515 = n8666 & n23514;
  assign n23516 = ~n7236 & n23515;
  assign n23517 = ~n6137 & n23516;
  assign n23518 = n6193 & n23517;
  assign n23519 = n6134 & n23518;
  assign n23520 = ~n7235 & n23519;
  assign n23521 = n7296 & n23520;
  assign n23522 = n7231 & n23521;
  assign n23523 = ~n23501 & ~n23522;
  assign n23524 = ~n23498 & n23523;
  assign n23525 = ~n23494 & n23524;
  assign n23526 = pi153 & ~n7663;
  assign n23527 = n8360 & n23526;
  assign n23528 = n8368 & n23527;
  assign n23529 = ~n7869 & n23528;
  assign n23530 = ~n8017 & n23529;
  assign n23531 = ~n8045 & n23530;
  assign n23532 = ~n8335 & n23531;
  assign n23533 = n8331 & n23532;
  assign n23534 = n8328 & n23533;
  assign n23535 = n8306 & n23534;
  assign n23536 = n8193 & n22073;
  assign n23537 = ~n5808 & n23536;
  assign n23538 = ~n6056 & n23537;
  assign n23539 = ~n8161 & n23538;
  assign n23540 = ~n8017 & n23539;
  assign n23541 = ~n7073 & n23540;
  assign n23542 = ~n8160 & n23541;
  assign n23543 = n8176 & n23542;
  assign n23544 = n8159 & n23543;
  assign n23545 = n8154 & n23544;
  assign n23546 = ~n23535 & ~n23545;
  assign n23547 = n23525 & n23546;
  assign n23548 = n23482 & n23547;
  assign n23549 = pi161 & ~n8391;
  assign n23550 = ~po161 & n23549;
  assign n23551 = ~n8017 & n23550;
  assign n23552 = ~n8314 & n23551;
  assign n23553 = n8281 & n23552;
  assign n23554 = n8390 & n23553;
  assign n23555 = n8383 & n23554;
  assign n23556 = n8264 & n22046;
  assign n23557 = ~n6784 & n23556;
  assign n23558 = ~n8232 & n23557;
  assign n23559 = ~n8017 & n23558;
  assign n23560 = ~n7158 & n23559;
  assign n23561 = ~n8231 & n23560;
  assign n23562 = n8247 & n23561;
  assign n23563 = n8230 & n23562;
  assign n23564 = n8227 & n23563;
  assign n23565 = pi145 & ~n6754;
  assign n23566 = ~n8017 & n23565;
  assign n23567 = ~n7204 & n23566;
  assign n23568 = ~n8282 & n23567;
  assign n23569 = n8288 & n23568;
  assign n23570 = n8281 & n23569;
  assign n23571 = n8280 & n23570;
  assign n23572 = ~n23564 & ~n23571;
  assign n23573 = ~n23555 & n23572;
  assign n23574 = ~n1958 & n18933;
  assign n23575 = n7910 & n23574;
  assign n23576 = ~n2242 & n23575;
  assign n23577 = ~n3095 & n23576;
  assign n23578 = ~n3997 & n23577;
  assign n23579 = ~n4003 & n23578;
  assign n23580 = ~n4837 & n23579;
  assign n23581 = ~n5822 & n23580;
  assign n23582 = ~n6820 & n23581;
  assign n23583 = ~n7907 & n23582;
  assign n23584 = ~n7906 & n23583;
  assign n23585 = ~n7785 & n23584;
  assign n23586 = ~n7905 & n23585;
  assign n23587 = n7925 & n23586;
  assign n23588 = n7904 & n23587;
  assign n23589 = n7897 & n23588;
  assign n23590 = n7978 & n22056;
  assign n23591 = ~n3066 & n23590;
  assign n23592 = ~n3983 & n23591;
  assign n23593 = ~n4003 & n23592;
  assign n23594 = ~n4024 & n23593;
  assign n23595 = ~n4999 & n23594;
  assign n23596 = ~n5827 & n23595;
  assign n23597 = ~n7870 & n23596;
  assign n23598 = ~n7842 & n23597;
  assign n23599 = ~n6893 & n23598;
  assign n23600 = ~n7841 & n23599;
  assign n23601 = n7887 & n23600;
  assign n23602 = n7840 & n23601;
  assign n23603 = n7810 & n23602;
  assign n23604 = ~n23589 & ~n23603;
  assign n23605 = n8121 & n22119;
  assign n23606 = ~n4817 & n23605;
  assign n23607 = ~n4902 & n23606;
  assign n23608 = ~n6001 & n23607;
  assign n23609 = ~n8094 & n23608;
  assign n23610 = ~n8017 & n23609;
  assign n23611 = ~n7014 & n23610;
  assign n23612 = ~n8093 & n23611;
  assign n23613 = n8111 & n23612;
  assign n23614 = n8092 & n23613;
  assign n23615 = n8086 & n23614;
  assign n23616 = pi041 & ~n1115;
  assign n23617 = ~n1026 & n23616;
  assign n23618 = ~n1086 & n23617;
  assign n23619 = n1239 & n23618;
  assign n23620 = ~n1270 & n23619;
  assign n23621 = n844 & n23620;
  assign n23622 = ~n1372 & n23621;
  assign n23623 = ~n2243 & n23622;
  assign n23624 = ~n3104 & n23623;
  assign n23625 = ~n3971 & n23624;
  assign n23626 = ~n4003 & n23625;
  assign n23627 = ~n4872 & n23626;
  assign n23628 = ~n5801 & n23627;
  assign n23629 = ~n6739 & n23628;
  assign n23630 = ~n7945 & n23629;
  assign n23631 = ~n7944 & n23630;
  assign n23632 = ~n7807 & n23631;
  assign n23633 = ~n7943 & n23632;
  assign n23634 = n7966 & n23633;
  assign n23635 = n7942 & n23634;
  assign n23636 = n7935 & n23635;
  assign n23637 = ~n23615 & ~n23636;
  assign n23638 = n23604 & n23637;
  assign n23639 = n23573 & n23638;
  assign po090 = ~n23548 | ~n23639;
  assign n23641 = ~n6967 & n22343;
  assign n23642 = ~n8017 & n23641;
  assign n23643 = ~n8044 & n23642;
  assign n23644 = n8052 & n23643;
  assign n23645 = ~n6114 & n21182;
  assign n23646 = ~n7095 & n23645;
  assign n23647 = ~n8017 & n23646;
  assign n23648 = n8155 & n23647;
  assign n23649 = n8216 & n23648;
  assign n23650 = n8210 & n23649;
  assign n23651 = ~n7029 & n22316;
  assign n23652 = ~n8017 & n23651;
  assign n23653 = ~n8045 & n23652;
  assign n23654 = n8143 & n23653;
  assign n23655 = n8137 & n23654;
  assign n23656 = ~n23650 & ~n23655;
  assign n23657 = ~n23644 & n23656;
  assign n23658 = n8059 & n22244;
  assign n23659 = ~n3940 & n23658;
  assign n23660 = ~n4001 & n23659;
  assign n23661 = ~n5043 & n23660;
  assign n23662 = ~n5943 & n23661;
  assign n23663 = ~n8018 & n23662;
  assign n23664 = ~n8017 & n23663;
  assign n23665 = ~n6951 & n23664;
  assign n23666 = ~n8016 & n23665;
  assign n23667 = n8034 & n23666;
  assign n23668 = n8015 & n23667;
  assign n23669 = n8008 & n23668;
  assign n23670 = pi178 & ~n501;
  assign n23671 = n5714 & n23670;
  assign n23672 = n5719 & n23671;
  assign n23673 = n8912 & n23672;
  assign n23674 = ~n1172 & n23673;
  assign n23675 = ~n996 & n23674;
  assign n23676 = ~n2306 & n23675;
  assign n23677 = ~n500 & n23676;
  assign n23678 = n6677 & n23677;
  assign n23679 = n8880 & n23678;
  assign n23680 = n7284 & n23679;
  assign n23681 = ~n7236 & n23680;
  assign n23682 = ~n6137 & n23681;
  assign n23683 = n6193 & n23682;
  assign n23684 = n6134 & n23683;
  assign n23685 = ~n8867 & n23684;
  assign n23686 = ~n7235 & n23685;
  assign n23687 = n7296 & n23686;
  assign n23688 = n7231 & n23687;
  assign n23689 = ~n8866 & n23688;
  assign n23690 = n8898 & n23689;
  assign n23691 = n8863 & n23690;
  assign n23692 = ~n6917 & n22347;
  assign n23693 = ~n7993 & n23692;
  assign n23694 = n7998 & n23693;
  assign n23695 = pi170 & ~n501;
  assign n23696 = n8692 & n23695;
  assign n23697 = n8941 & n23696;
  assign n23698 = n8946 & n23697;
  assign n23699 = n8940 & n23698;
  assign n23700 = ~n1172 & n23699;
  assign n23701 = ~n1025 & n23700;
  assign n23702 = ~n996 & n23701;
  assign n23703 = n8701 & n23702;
  assign n23704 = n3821 & n23703;
  assign n23705 = n8681 & n23704;
  assign n23706 = n8824 & n23705;
  assign n23707 = n8679 & n23706;
  assign n23708 = n8666 & n23707;
  assign n23709 = ~n7236 & n23708;
  assign n23710 = ~n6137 & n23709;
  assign n23711 = n6193 & n23710;
  assign n23712 = n6134 & n23711;
  assign n23713 = ~n7235 & n23712;
  assign n23714 = n7296 & n23713;
  assign n23715 = n7231 & n23714;
  assign n23716 = ~n23694 & ~n23715;
  assign n23717 = ~n23691 & n23716;
  assign n23718 = ~n23669 & n23717;
  assign n23719 = pi042 & ~n1115;
  assign n23720 = ~n1026 & n23719;
  assign n23721 = ~n1086 & n23720;
  assign n23722 = n1239 & n23721;
  assign n23723 = ~n1270 & n23722;
  assign n23724 = n844 & n23723;
  assign n23725 = ~n1372 & n23724;
  assign n23726 = ~n2243 & n23725;
  assign n23727 = ~n3104 & n23726;
  assign n23728 = ~n3971 & n23727;
  assign n23729 = ~n4003 & n23728;
  assign n23730 = ~n4872 & n23729;
  assign n23731 = ~n5801 & n23730;
  assign n23732 = ~n6739 & n23731;
  assign n23733 = ~n7945 & n23732;
  assign n23734 = ~n7944 & n23733;
  assign n23735 = ~n7807 & n23734;
  assign n23736 = ~n7943 & n23735;
  assign n23737 = n7966 & n23736;
  assign n23738 = n7942 & n23737;
  assign n23739 = n7935 & n23738;
  assign n23740 = n8264 & n22271;
  assign n23741 = ~n6784 & n23740;
  assign n23742 = ~n8232 & n23741;
  assign n23743 = ~n8017 & n23742;
  assign n23744 = ~n7158 & n23743;
  assign n23745 = ~n8231 & n23744;
  assign n23746 = n8247 & n23745;
  assign n23747 = n8230 & n23746;
  assign n23748 = n8227 & n23747;
  assign n23749 = ~n23739 & ~n23748;
  assign n23750 = n23718 & n23749;
  assign n23751 = n23657 & n23750;
  assign n23752 = pi154 & ~n7663;
  assign n23753 = n8360 & n23752;
  assign n23754 = n8368 & n23753;
  assign n23755 = ~n7869 & n23754;
  assign n23756 = ~n8017 & n23755;
  assign n23757 = ~n8045 & n23756;
  assign n23758 = ~n8335 & n23757;
  assign n23759 = n8331 & n23758;
  assign n23760 = n8328 & n23759;
  assign n23761 = n8306 & n23760;
  assign n23762 = pi162 & ~n8391;
  assign n23763 = ~po161 & n23762;
  assign n23764 = ~n8017 & n23763;
  assign n23765 = ~n8314 & n23764;
  assign n23766 = n8281 & n23765;
  assign n23767 = n8390 & n23766;
  assign n23768 = n8383 & n23767;
  assign n23769 = n8193 & n22231;
  assign n23770 = ~n5808 & n23769;
  assign n23771 = ~n6056 & n23770;
  assign n23772 = ~n8161 & n23771;
  assign n23773 = ~n8017 & n23772;
  assign n23774 = ~n7073 & n23773;
  assign n23775 = ~n8160 & n23774;
  assign n23776 = n8176 & n23775;
  assign n23777 = n8159 & n23776;
  assign n23778 = n8154 & n23777;
  assign n23779 = ~n23768 & ~n23778;
  assign n23780 = ~n23761 & n23779;
  assign n23781 = pi146 & ~n6754;
  assign n23782 = ~n8017 & n23781;
  assign n23783 = ~n7204 & n23782;
  assign n23784 = ~n8282 & n23783;
  assign n23785 = n8288 & n23784;
  assign n23786 = n8281 & n23785;
  assign n23787 = n8280 & n23786;
  assign n23788 = ~n1958 & n18992;
  assign n23789 = n7910 & n23788;
  assign n23790 = ~n2242 & n23789;
  assign n23791 = ~n3095 & n23790;
  assign n23792 = ~n3997 & n23791;
  assign n23793 = ~n4003 & n23792;
  assign n23794 = ~n4837 & n23793;
  assign n23795 = ~n5822 & n23794;
  assign n23796 = ~n6820 & n23795;
  assign n23797 = ~n7907 & n23796;
  assign n23798 = ~n7906 & n23797;
  assign n23799 = ~n7785 & n23798;
  assign n23800 = ~n7905 & n23799;
  assign n23801 = n7925 & n23800;
  assign n23802 = n7904 & n23801;
  assign n23803 = n7897 & n23802;
  assign n23804 = ~n23787 & ~n23803;
  assign n23805 = n7978 & n22281;
  assign n23806 = ~n3066 & n23805;
  assign n23807 = ~n3983 & n23806;
  assign n23808 = ~n4003 & n23807;
  assign n23809 = ~n4024 & n23808;
  assign n23810 = ~n4999 & n23809;
  assign n23811 = ~n5827 & n23810;
  assign n23812 = ~n7870 & n23811;
  assign n23813 = ~n7842 & n23812;
  assign n23814 = ~n6893 & n23813;
  assign n23815 = ~n7841 & n23814;
  assign n23816 = n7887 & n23815;
  assign n23817 = n7840 & n23816;
  assign n23818 = n7810 & n23817;
  assign n23819 = n8121 & n22257;
  assign n23820 = ~n4817 & n23819;
  assign n23821 = ~n4902 & n23820;
  assign n23822 = ~n6001 & n23821;
  assign n23823 = ~n8094 & n23822;
  assign n23824 = ~n8017 & n23823;
  assign n23825 = ~n7014 & n23824;
  assign n23826 = ~n8093 & n23825;
  assign n23827 = n8111 & n23826;
  assign n23828 = n8092 & n23827;
  assign n23829 = n8086 & n23828;
  assign n23830 = ~n23818 & ~n23829;
  assign n23831 = n23804 & n23830;
  assign n23832 = n23780 & n23831;
  assign po091 = ~n23751 | ~n23832;
  assign n23834 = ~n6967 & n22510;
  assign n23835 = ~n8017 & n23834;
  assign n23836 = ~n8044 & n23835;
  assign n23837 = n8052 & n23836;
  assign n23838 = ~n6114 & n21308;
  assign n23839 = ~n7095 & n23838;
  assign n23840 = ~n8017 & n23839;
  assign n23841 = n8155 & n23840;
  assign n23842 = n8216 & n23841;
  assign n23843 = n8210 & n23842;
  assign n23844 = ~n7029 & n22483;
  assign n23845 = ~n8017 & n23844;
  assign n23846 = ~n8045 & n23845;
  assign n23847 = n8143 & n23846;
  assign n23848 = n8137 & n23847;
  assign n23849 = ~n23843 & ~n23848;
  assign n23850 = ~n23837 & n23849;
  assign n23851 = pi043 & ~n1115;
  assign n23852 = ~n1026 & n23851;
  assign n23853 = ~n1086 & n23852;
  assign n23854 = n1239 & n23853;
  assign n23855 = ~n1270 & n23854;
  assign n23856 = n844 & n23855;
  assign n23857 = ~n1372 & n23856;
  assign n23858 = ~n2243 & n23857;
  assign n23859 = ~n3104 & n23858;
  assign n23860 = ~n3971 & n23859;
  assign n23861 = ~n4003 & n23860;
  assign n23862 = ~n4872 & n23861;
  assign n23863 = ~n5801 & n23862;
  assign n23864 = ~n6739 & n23863;
  assign n23865 = ~n7945 & n23864;
  assign n23866 = ~n7944 & n23865;
  assign n23867 = ~n7807 & n23866;
  assign n23868 = ~n7943 & n23867;
  assign n23869 = n7966 & n23868;
  assign n23870 = n7942 & n23869;
  assign n23871 = n7935 & n23870;
  assign n23872 = pi179 & ~n501;
  assign n23873 = n5714 & n23872;
  assign n23874 = n5719 & n23873;
  assign n23875 = n8912 & n23874;
  assign n23876 = ~n1172 & n23875;
  assign n23877 = ~n996 & n23876;
  assign n23878 = ~n2306 & n23877;
  assign n23879 = ~n500 & n23878;
  assign n23880 = n6677 & n23879;
  assign n23881 = n8880 & n23880;
  assign n23882 = n7284 & n23881;
  assign n23883 = ~n7236 & n23882;
  assign n23884 = ~n6137 & n23883;
  assign n23885 = n6193 & n23884;
  assign n23886 = n6134 & n23885;
  assign n23887 = ~n8867 & n23886;
  assign n23888 = ~n7235 & n23887;
  assign n23889 = n7296 & n23888;
  assign n23890 = n7231 & n23889;
  assign n23891 = ~n8866 & n23890;
  assign n23892 = n8898 & n23891;
  assign n23893 = n8863 & n23892;
  assign n23894 = ~n6917 & n22514;
  assign n23895 = ~n7993 & n23894;
  assign n23896 = n7998 & n23895;
  assign n23897 = pi171 & ~n501;
  assign n23898 = n8692 & n23897;
  assign n23899 = n8941 & n23898;
  assign n23900 = n8946 & n23899;
  assign n23901 = n8940 & n23900;
  assign n23902 = ~n1172 & n23901;
  assign n23903 = ~n1025 & n23902;
  assign n23904 = ~n996 & n23903;
  assign n23905 = n8701 & n23904;
  assign n23906 = n3821 & n23905;
  assign n23907 = n8681 & n23906;
  assign n23908 = n8824 & n23907;
  assign n23909 = n8679 & n23908;
  assign n23910 = n8666 & n23909;
  assign n23911 = ~n7236 & n23910;
  assign n23912 = ~n6137 & n23911;
  assign n23913 = n6193 & n23912;
  assign n23914 = n6134 & n23913;
  assign n23915 = ~n7235 & n23914;
  assign n23916 = n7296 & n23915;
  assign n23917 = n7231 & n23916;
  assign n23918 = ~n23896 & ~n23917;
  assign n23919 = ~n23893 & n23918;
  assign n23920 = ~n23871 & n23919;
  assign n23921 = n8264 & n22438;
  assign n23922 = ~n6784 & n23921;
  assign n23923 = ~n8232 & n23922;
  assign n23924 = ~n8017 & n23923;
  assign n23925 = ~n7158 & n23924;
  assign n23926 = ~n8231 & n23925;
  assign n23927 = n8247 & n23926;
  assign n23928 = n8230 & n23927;
  assign n23929 = n8227 & n23928;
  assign n23930 = n8059 & n22411;
  assign n23931 = ~n3940 & n23930;
  assign n23932 = ~n4001 & n23931;
  assign n23933 = ~n5043 & n23932;
  assign n23934 = ~n5943 & n23933;
  assign n23935 = ~n8018 & n23934;
  assign n23936 = ~n8017 & n23935;
  assign n23937 = ~n6951 & n23936;
  assign n23938 = ~n8016 & n23937;
  assign n23939 = n8034 & n23938;
  assign n23940 = n8015 & n23939;
  assign n23941 = n8008 & n23940;
  assign n23942 = ~n23929 & ~n23941;
  assign n23943 = n23920 & n23942;
  assign n23944 = n23850 & n23943;
  assign n23945 = pi155 & ~n7663;
  assign n23946 = n8360 & n23945;
  assign n23947 = n8368 & n23946;
  assign n23948 = ~n7869 & n23947;
  assign n23949 = ~n8017 & n23948;
  assign n23950 = ~n8045 & n23949;
  assign n23951 = ~n8335 & n23950;
  assign n23952 = n8331 & n23951;
  assign n23953 = n8328 & n23952;
  assign n23954 = n8306 & n23953;
  assign n23955 = pi163 & ~n8391;
  assign n23956 = ~po161 & n23955;
  assign n23957 = ~n8017 & n23956;
  assign n23958 = ~n8314 & n23957;
  assign n23959 = n8281 & n23958;
  assign n23960 = n8390 & n23959;
  assign n23961 = n8383 & n23960;
  assign n23962 = n8193 & n22398;
  assign n23963 = ~n5808 & n23962;
  assign n23964 = ~n6056 & n23963;
  assign n23965 = ~n8161 & n23964;
  assign n23966 = ~n8017 & n23965;
  assign n23967 = ~n7073 & n23966;
  assign n23968 = ~n8160 & n23967;
  assign n23969 = n8176 & n23968;
  assign n23970 = n8159 & n23969;
  assign n23971 = n8154 & n23970;
  assign n23972 = ~n23961 & ~n23971;
  assign n23973 = ~n23954 & n23972;
  assign n23974 = n7978 & n22448;
  assign n23975 = ~n3066 & n23974;
  assign n23976 = ~n3983 & n23975;
  assign n23977 = ~n4003 & n23976;
  assign n23978 = ~n4024 & n23977;
  assign n23979 = ~n4999 & n23978;
  assign n23980 = ~n5827 & n23979;
  assign n23981 = ~n7870 & n23980;
  assign n23982 = ~n7842 & n23981;
  assign n23983 = ~n6893 & n23982;
  assign n23984 = ~n7841 & n23983;
  assign n23985 = n7887 & n23984;
  assign n23986 = n7840 & n23985;
  assign n23987 = n7810 & n23986;
  assign n23988 = pi147 & ~n6754;
  assign n23989 = ~n8017 & n23988;
  assign n23990 = ~n7204 & n23989;
  assign n23991 = ~n8282 & n23990;
  assign n23992 = n8288 & n23991;
  assign n23993 = n8281 & n23992;
  assign n23994 = n8280 & n23993;
  assign n23995 = ~n23987 & ~n23994;
  assign n23996 = ~n1958 & n19051;
  assign n23997 = n7910 & n23996;
  assign n23998 = ~n2242 & n23997;
  assign n23999 = ~n3095 & n23998;
  assign n24000 = ~n3997 & n23999;
  assign n24001 = ~n4003 & n24000;
  assign n24002 = ~n4837 & n24001;
  assign n24003 = ~n5822 & n24002;
  assign n24004 = ~n6820 & n24003;
  assign n24005 = ~n7907 & n24004;
  assign n24006 = ~n7906 & n24005;
  assign n24007 = ~n7785 & n24006;
  assign n24008 = ~n7905 & n24007;
  assign n24009 = n7925 & n24008;
  assign n24010 = n7904 & n24009;
  assign n24011 = n7897 & n24010;
  assign n24012 = n8121 & n22424;
  assign n24013 = ~n4817 & n24012;
  assign n24014 = ~n4902 & n24013;
  assign n24015 = ~n6001 & n24014;
  assign n24016 = ~n8094 & n24015;
  assign n24017 = ~n8017 & n24016;
  assign n24018 = ~n7014 & n24017;
  assign n24019 = ~n8093 & n24018;
  assign n24020 = n8111 & n24019;
  assign n24021 = n8092 & n24020;
  assign n24022 = n8086 & n24021;
  assign n24023 = ~n24011 & ~n24022;
  assign n24024 = n23995 & n24023;
  assign n24025 = n23973 & n24024;
  assign po092 = ~n23944 | ~n24025;
  assign n24027 = pi180 & ~n501;
  assign n24028 = n5714 & n24027;
  assign n24029 = n5719 & n24028;
  assign n24030 = n8912 & n24029;
  assign n24031 = ~n1172 & n24030;
  assign n24032 = ~n996 & n24031;
  assign n24033 = ~n2306 & n24032;
  assign n24034 = ~n500 & n24033;
  assign n24035 = n6677 & n24034;
  assign n24036 = n8880 & n24035;
  assign n24037 = n7284 & n24036;
  assign n24038 = ~n7236 & n24037;
  assign n24039 = ~n6137 & n24038;
  assign n24040 = n6193 & n24039;
  assign n24041 = n6134 & n24040;
  assign n24042 = ~n8867 & n24041;
  assign n24043 = ~n7235 & n24042;
  assign n24044 = n7296 & n24043;
  assign n24045 = n7231 & n24044;
  assign n24046 = ~n8866 & n24045;
  assign n24047 = n8898 & n24046;
  assign n24048 = n8863 & n24047;
  assign n24049 = ~n7029 & n22650;
  assign n24050 = ~n8017 & n24049;
  assign n24051 = ~n8045 & n24050;
  assign n24052 = n8143 & n24051;
  assign n24053 = n8137 & n24052;
  assign n24054 = ~n6967 & n22677;
  assign n24055 = ~n8017 & n24054;
  assign n24056 = ~n8044 & n24055;
  assign n24057 = n8052 & n24056;
  assign n24058 = ~n24053 & ~n24057;
  assign n24059 = ~n24048 & n24058;
  assign n24060 = n8059 & n22578;
  assign n24061 = ~n3940 & n24060;
  assign n24062 = ~n4001 & n24061;
  assign n24063 = ~n5043 & n24062;
  assign n24064 = ~n5943 & n24063;
  assign n24065 = ~n8018 & n24064;
  assign n24066 = ~n8017 & n24065;
  assign n24067 = ~n6951 & n24066;
  assign n24068 = ~n8016 & n24067;
  assign n24069 = n8034 & n24068;
  assign n24070 = n8015 & n24069;
  assign n24071 = n8008 & n24070;
  assign n24072 = ~n6114 & n21434;
  assign n24073 = ~n7095 & n24072;
  assign n24074 = ~n8017 & n24073;
  assign n24075 = n8155 & n24074;
  assign n24076 = n8216 & n24075;
  assign n24077 = n8210 & n24076;
  assign n24078 = ~n6917 & n22681;
  assign n24079 = ~n7993 & n24078;
  assign n24080 = n7998 & n24079;
  assign n24081 = pi172 & ~n501;
  assign n24082 = n8692 & n24081;
  assign n24083 = n8941 & n24082;
  assign n24084 = n8946 & n24083;
  assign n24085 = n8940 & n24084;
  assign n24086 = ~n1172 & n24085;
  assign n24087 = ~n1025 & n24086;
  assign n24088 = ~n996 & n24087;
  assign n24089 = n8701 & n24088;
  assign n24090 = n3821 & n24089;
  assign n24091 = n8681 & n24090;
  assign n24092 = n8824 & n24091;
  assign n24093 = n8679 & n24092;
  assign n24094 = n8666 & n24093;
  assign n24095 = ~n7236 & n24094;
  assign n24096 = ~n6137 & n24095;
  assign n24097 = n6193 & n24096;
  assign n24098 = n6134 & n24097;
  assign n24099 = ~n7235 & n24098;
  assign n24100 = n7296 & n24099;
  assign n24101 = n7231 & n24100;
  assign n24102 = ~n24080 & ~n24101;
  assign n24103 = ~n24077 & n24102;
  assign n24104 = ~n24071 & n24103;
  assign n24105 = pi044 & ~n1115;
  assign n24106 = ~n1026 & n24105;
  assign n24107 = ~n1086 & n24106;
  assign n24108 = n1239 & n24107;
  assign n24109 = ~n1270 & n24108;
  assign n24110 = n844 & n24109;
  assign n24111 = ~n1372 & n24110;
  assign n24112 = ~n2243 & n24111;
  assign n24113 = ~n3104 & n24112;
  assign n24114 = ~n3971 & n24113;
  assign n24115 = ~n4003 & n24114;
  assign n24116 = ~n4872 & n24115;
  assign n24117 = ~n5801 & n24116;
  assign n24118 = ~n6739 & n24117;
  assign n24119 = ~n7945 & n24118;
  assign n24120 = ~n7944 & n24119;
  assign n24121 = ~n7807 & n24120;
  assign n24122 = ~n7943 & n24121;
  assign n24123 = n7966 & n24122;
  assign n24124 = n7942 & n24123;
  assign n24125 = n7935 & n24124;
  assign n24126 = n8264 & n22605;
  assign n24127 = ~n6784 & n24126;
  assign n24128 = ~n8232 & n24127;
  assign n24129 = ~n8017 & n24128;
  assign n24130 = ~n7158 & n24129;
  assign n24131 = ~n8231 & n24130;
  assign n24132 = n8247 & n24131;
  assign n24133 = n8230 & n24132;
  assign n24134 = n8227 & n24133;
  assign n24135 = ~n24125 & ~n24134;
  assign n24136 = n24104 & n24135;
  assign n24137 = n24059 & n24136;
  assign n24138 = ~n1958 & n19110;
  assign n24139 = n7910 & n24138;
  assign n24140 = ~n2242 & n24139;
  assign n24141 = ~n3095 & n24140;
  assign n24142 = ~n3997 & n24141;
  assign n24143 = ~n4003 & n24142;
  assign n24144 = ~n4837 & n24143;
  assign n24145 = ~n5822 & n24144;
  assign n24146 = ~n6820 & n24145;
  assign n24147 = ~n7907 & n24146;
  assign n24148 = ~n7906 & n24147;
  assign n24149 = ~n7785 & n24148;
  assign n24150 = ~n7905 & n24149;
  assign n24151 = n7925 & n24150;
  assign n24152 = n7904 & n24151;
  assign n24153 = n7897 & n24152;
  assign n24154 = n7978 & n22615;
  assign n24155 = ~n3066 & n24154;
  assign n24156 = ~n3983 & n24155;
  assign n24157 = ~n4003 & n24156;
  assign n24158 = ~n4024 & n24157;
  assign n24159 = ~n4999 & n24158;
  assign n24160 = ~n5827 & n24159;
  assign n24161 = ~n7870 & n24160;
  assign n24162 = ~n7842 & n24161;
  assign n24163 = ~n6893 & n24162;
  assign n24164 = ~n7841 & n24163;
  assign n24165 = n7887 & n24164;
  assign n24166 = n7840 & n24165;
  assign n24167 = n7810 & n24166;
  assign n24168 = pi148 & ~n6754;
  assign n24169 = ~n8017 & n24168;
  assign n24170 = ~n7204 & n24169;
  assign n24171 = ~n8282 & n24170;
  assign n24172 = n8288 & n24171;
  assign n24173 = n8281 & n24172;
  assign n24174 = n8280 & n24173;
  assign n24175 = ~n24167 & ~n24174;
  assign n24176 = ~n24153 & n24175;
  assign n24177 = n8121 & n22591;
  assign n24178 = ~n4817 & n24177;
  assign n24179 = ~n4902 & n24178;
  assign n24180 = ~n6001 & n24179;
  assign n24181 = ~n8094 & n24180;
  assign n24182 = ~n8017 & n24181;
  assign n24183 = ~n7014 & n24182;
  assign n24184 = ~n8093 & n24183;
  assign n24185 = n8111 & n24184;
  assign n24186 = n8092 & n24185;
  assign n24187 = n8086 & n24186;
  assign n24188 = pi164 & ~n8391;
  assign n24189 = ~po161 & n24188;
  assign n24190 = ~n8017 & n24189;
  assign n24191 = ~n8314 & n24190;
  assign n24192 = n8281 & n24191;
  assign n24193 = n8390 & n24192;
  assign n24194 = n8383 & n24193;
  assign n24195 = ~n24187 & ~n24194;
  assign n24196 = n8193 & n22565;
  assign n24197 = ~n5808 & n24196;
  assign n24198 = ~n6056 & n24197;
  assign n24199 = ~n8161 & n24198;
  assign n24200 = ~n8017 & n24199;
  assign n24201 = ~n7073 & n24200;
  assign n24202 = ~n8160 & n24201;
  assign n24203 = n8176 & n24202;
  assign n24204 = n8159 & n24203;
  assign n24205 = n8154 & n24204;
  assign n24206 = pi156 & ~n7663;
  assign n24207 = n8360 & n24206;
  assign n24208 = n8368 & n24207;
  assign n24209 = ~n7869 & n24208;
  assign n24210 = ~n8017 & n24209;
  assign n24211 = ~n8045 & n24210;
  assign n24212 = ~n8335 & n24211;
  assign n24213 = n8331 & n24212;
  assign n24214 = n8328 & n24213;
  assign n24215 = n8306 & n24214;
  assign n24216 = ~n24205 & ~n24215;
  assign n24217 = n24195 & n24216;
  assign n24218 = n24176 & n24217;
  assign po093 = ~n24137 | ~n24218;
  assign n24220 = pi181 & ~n501;
  assign n24221 = n5714 & n24220;
  assign n24222 = n5719 & n24221;
  assign n24223 = n8912 & n24222;
  assign n24224 = ~n1172 & n24223;
  assign n24225 = ~n996 & n24224;
  assign n24226 = ~n2306 & n24225;
  assign n24227 = ~n500 & n24226;
  assign n24228 = n6677 & n24227;
  assign n24229 = n8880 & n24228;
  assign n24230 = n7284 & n24229;
  assign n24231 = ~n7236 & n24230;
  assign n24232 = ~n6137 & n24231;
  assign n24233 = n6193 & n24232;
  assign n24234 = n6134 & n24233;
  assign n24235 = ~n8867 & n24234;
  assign n24236 = ~n7235 & n24235;
  assign n24237 = n7296 & n24236;
  assign n24238 = n7231 & n24237;
  assign n24239 = ~n8866 & n24238;
  assign n24240 = n8898 & n24239;
  assign n24241 = n8863 & n24240;
  assign n24242 = ~n7029 & n22817;
  assign n24243 = ~n8017 & n24242;
  assign n24244 = ~n8045 & n24243;
  assign n24245 = n8143 & n24244;
  assign n24246 = n8137 & n24245;
  assign n24247 = ~n6967 & n22844;
  assign n24248 = ~n8017 & n24247;
  assign n24249 = ~n8044 & n24248;
  assign n24250 = n8052 & n24249;
  assign n24251 = ~n24246 & ~n24250;
  assign n24252 = ~n24241 & n24251;
  assign n24253 = n8059 & n22745;
  assign n24254 = ~n3940 & n24253;
  assign n24255 = ~n4001 & n24254;
  assign n24256 = ~n5043 & n24255;
  assign n24257 = ~n5943 & n24256;
  assign n24258 = ~n8018 & n24257;
  assign n24259 = ~n8017 & n24258;
  assign n24260 = ~n6951 & n24259;
  assign n24261 = ~n8016 & n24260;
  assign n24262 = n8034 & n24261;
  assign n24263 = n8015 & n24262;
  assign n24264 = n8008 & n24263;
  assign n24265 = ~n6114 & n21560;
  assign n24266 = ~n7095 & n24265;
  assign n24267 = ~n8017 & n24266;
  assign n24268 = n8155 & n24267;
  assign n24269 = n8216 & n24268;
  assign n24270 = n8210 & n24269;
  assign n24271 = ~n6917 & n22848;
  assign n24272 = ~n7993 & n24271;
  assign n24273 = n7998 & n24272;
  assign n24274 = pi173 & ~n501;
  assign n24275 = n8692 & n24274;
  assign n24276 = n8941 & n24275;
  assign n24277 = n8946 & n24276;
  assign n24278 = n8940 & n24277;
  assign n24279 = ~n1172 & n24278;
  assign n24280 = ~n1025 & n24279;
  assign n24281 = ~n996 & n24280;
  assign n24282 = n8701 & n24281;
  assign n24283 = n3821 & n24282;
  assign n24284 = n8681 & n24283;
  assign n24285 = n8824 & n24284;
  assign n24286 = n8679 & n24285;
  assign n24287 = n8666 & n24286;
  assign n24288 = ~n7236 & n24287;
  assign n24289 = ~n6137 & n24288;
  assign n24290 = n6193 & n24289;
  assign n24291 = n6134 & n24290;
  assign n24292 = ~n7235 & n24291;
  assign n24293 = n7296 & n24292;
  assign n24294 = n7231 & n24293;
  assign n24295 = ~n24273 & ~n24294;
  assign n24296 = ~n24270 & n24295;
  assign n24297 = ~n24264 & n24296;
  assign n24298 = pi045 & ~n1115;
  assign n24299 = ~n1026 & n24298;
  assign n24300 = ~n1086 & n24299;
  assign n24301 = n1239 & n24300;
  assign n24302 = ~n1270 & n24301;
  assign n24303 = n844 & n24302;
  assign n24304 = ~n1372 & n24303;
  assign n24305 = ~n2243 & n24304;
  assign n24306 = ~n3104 & n24305;
  assign n24307 = ~n3971 & n24306;
  assign n24308 = ~n4003 & n24307;
  assign n24309 = ~n4872 & n24308;
  assign n24310 = ~n5801 & n24309;
  assign n24311 = ~n6739 & n24310;
  assign n24312 = ~n7945 & n24311;
  assign n24313 = ~n7944 & n24312;
  assign n24314 = ~n7807 & n24313;
  assign n24315 = ~n7943 & n24314;
  assign n24316 = n7966 & n24315;
  assign n24317 = n7942 & n24316;
  assign n24318 = n7935 & n24317;
  assign n24319 = n8264 & n22772;
  assign n24320 = ~n6784 & n24319;
  assign n24321 = ~n8232 & n24320;
  assign n24322 = ~n8017 & n24321;
  assign n24323 = ~n7158 & n24322;
  assign n24324 = ~n8231 & n24323;
  assign n24325 = n8247 & n24324;
  assign n24326 = n8230 & n24325;
  assign n24327 = n8227 & n24326;
  assign n24328 = ~n24318 & ~n24327;
  assign n24329 = n24297 & n24328;
  assign n24330 = n24252 & n24329;
  assign n24331 = ~n1958 & n19169;
  assign n24332 = n7910 & n24331;
  assign n24333 = ~n2242 & n24332;
  assign n24334 = ~n3095 & n24333;
  assign n24335 = ~n3997 & n24334;
  assign n24336 = ~n4003 & n24335;
  assign n24337 = ~n4837 & n24336;
  assign n24338 = ~n5822 & n24337;
  assign n24339 = ~n6820 & n24338;
  assign n24340 = ~n7907 & n24339;
  assign n24341 = ~n7906 & n24340;
  assign n24342 = ~n7785 & n24341;
  assign n24343 = ~n7905 & n24342;
  assign n24344 = n7925 & n24343;
  assign n24345 = n7904 & n24344;
  assign n24346 = n7897 & n24345;
  assign n24347 = n7978 & n22782;
  assign n24348 = ~n3066 & n24347;
  assign n24349 = ~n3983 & n24348;
  assign n24350 = ~n4003 & n24349;
  assign n24351 = ~n4024 & n24350;
  assign n24352 = ~n4999 & n24351;
  assign n24353 = ~n5827 & n24352;
  assign n24354 = ~n7870 & n24353;
  assign n24355 = ~n7842 & n24354;
  assign n24356 = ~n6893 & n24355;
  assign n24357 = ~n7841 & n24356;
  assign n24358 = n7887 & n24357;
  assign n24359 = n7840 & n24358;
  assign n24360 = n7810 & n24359;
  assign n24361 = pi149 & ~n6754;
  assign n24362 = ~n8017 & n24361;
  assign n24363 = ~n7204 & n24362;
  assign n24364 = ~n8282 & n24363;
  assign n24365 = n8288 & n24364;
  assign n24366 = n8281 & n24365;
  assign n24367 = n8280 & n24366;
  assign n24368 = ~n24360 & ~n24367;
  assign n24369 = ~n24346 & n24368;
  assign n24370 = n8121 & n22758;
  assign n24371 = ~n4817 & n24370;
  assign n24372 = ~n4902 & n24371;
  assign n24373 = ~n6001 & n24372;
  assign n24374 = ~n8094 & n24373;
  assign n24375 = ~n8017 & n24374;
  assign n24376 = ~n7014 & n24375;
  assign n24377 = ~n8093 & n24376;
  assign n24378 = n8111 & n24377;
  assign n24379 = n8092 & n24378;
  assign n24380 = n8086 & n24379;
  assign n24381 = pi165 & ~n8391;
  assign n24382 = ~po161 & n24381;
  assign n24383 = ~n8017 & n24382;
  assign n24384 = ~n8314 & n24383;
  assign n24385 = n8281 & n24384;
  assign n24386 = n8390 & n24385;
  assign n24387 = n8383 & n24386;
  assign n24388 = ~n24380 & ~n24387;
  assign n24389 = n8193 & n22732;
  assign n24390 = ~n5808 & n24389;
  assign n24391 = ~n6056 & n24390;
  assign n24392 = ~n8161 & n24391;
  assign n24393 = ~n8017 & n24392;
  assign n24394 = ~n7073 & n24393;
  assign n24395 = ~n8160 & n24394;
  assign n24396 = n8176 & n24395;
  assign n24397 = n8159 & n24396;
  assign n24398 = n8154 & n24397;
  assign n24399 = pi157 & ~n7663;
  assign n24400 = n8360 & n24399;
  assign n24401 = n8368 & n24400;
  assign n24402 = ~n7869 & n24401;
  assign n24403 = ~n8017 & n24402;
  assign n24404 = ~n8045 & n24403;
  assign n24405 = ~n8335 & n24404;
  assign n24406 = n8331 & n24405;
  assign n24407 = n8328 & n24406;
  assign n24408 = n8306 & n24407;
  assign n24409 = ~n24398 & ~n24408;
  assign n24410 = n24388 & n24409;
  assign n24411 = n24369 & n24410;
  assign po094 = ~n24330 | ~n24411;
  assign n24413 = pi182 & ~n501;
  assign n24414 = n5714 & n24413;
  assign n24415 = n5719 & n24414;
  assign n24416 = n8912 & n24415;
  assign n24417 = ~n1172 & n24416;
  assign n24418 = ~n996 & n24417;
  assign n24419 = ~n2306 & n24418;
  assign n24420 = ~n500 & n24419;
  assign n24421 = n6677 & n24420;
  assign n24422 = n8880 & n24421;
  assign n24423 = n7284 & n24422;
  assign n24424 = ~n7236 & n24423;
  assign n24425 = ~n6137 & n24424;
  assign n24426 = n6193 & n24425;
  assign n24427 = n6134 & n24426;
  assign n24428 = ~n8867 & n24427;
  assign n24429 = ~n7235 & n24428;
  assign n24430 = n7296 & n24429;
  assign n24431 = n7231 & n24430;
  assign n24432 = ~n8866 & n24431;
  assign n24433 = n8898 & n24432;
  assign n24434 = n8863 & n24433;
  assign n24435 = ~n7029 & n22984;
  assign n24436 = ~n8017 & n24435;
  assign n24437 = ~n8045 & n24436;
  assign n24438 = n8143 & n24437;
  assign n24439 = n8137 & n24438;
  assign n24440 = ~n6967 & n23011;
  assign n24441 = ~n8017 & n24440;
  assign n24442 = ~n8044 & n24441;
  assign n24443 = n8052 & n24442;
  assign n24444 = ~n24439 & ~n24443;
  assign n24445 = ~n24434 & n24444;
  assign n24446 = n8059 & n22912;
  assign n24447 = ~n3940 & n24446;
  assign n24448 = ~n4001 & n24447;
  assign n24449 = ~n5043 & n24448;
  assign n24450 = ~n5943 & n24449;
  assign n24451 = ~n8018 & n24450;
  assign n24452 = ~n8017 & n24451;
  assign n24453 = ~n6951 & n24452;
  assign n24454 = ~n8016 & n24453;
  assign n24455 = n8034 & n24454;
  assign n24456 = n8015 & n24455;
  assign n24457 = n8008 & n24456;
  assign n24458 = ~n6114 & n21686;
  assign n24459 = ~n7095 & n24458;
  assign n24460 = ~n8017 & n24459;
  assign n24461 = n8155 & n24460;
  assign n24462 = n8216 & n24461;
  assign n24463 = n8210 & n24462;
  assign n24464 = ~n6917 & n23015;
  assign n24465 = ~n7993 & n24464;
  assign n24466 = n7998 & n24465;
  assign n24467 = pi174 & ~n501;
  assign n24468 = n8692 & n24467;
  assign n24469 = n8941 & n24468;
  assign n24470 = n8946 & n24469;
  assign n24471 = n8940 & n24470;
  assign n24472 = ~n1172 & n24471;
  assign n24473 = ~n1025 & n24472;
  assign n24474 = ~n996 & n24473;
  assign n24475 = n8701 & n24474;
  assign n24476 = n3821 & n24475;
  assign n24477 = n8681 & n24476;
  assign n24478 = n8824 & n24477;
  assign n24479 = n8679 & n24478;
  assign n24480 = n8666 & n24479;
  assign n24481 = ~n7236 & n24480;
  assign n24482 = ~n6137 & n24481;
  assign n24483 = n6193 & n24482;
  assign n24484 = n6134 & n24483;
  assign n24485 = ~n7235 & n24484;
  assign n24486 = n7296 & n24485;
  assign n24487 = n7231 & n24486;
  assign n24488 = ~n24466 & ~n24487;
  assign n24489 = ~n24463 & n24488;
  assign n24490 = ~n24457 & n24489;
  assign n24491 = pi046 & ~n1115;
  assign n24492 = ~n1026 & n24491;
  assign n24493 = ~n1086 & n24492;
  assign n24494 = n1239 & n24493;
  assign n24495 = ~n1270 & n24494;
  assign n24496 = n844 & n24495;
  assign n24497 = ~n1372 & n24496;
  assign n24498 = ~n2243 & n24497;
  assign n24499 = ~n3104 & n24498;
  assign n24500 = ~n3971 & n24499;
  assign n24501 = ~n4003 & n24500;
  assign n24502 = ~n4872 & n24501;
  assign n24503 = ~n5801 & n24502;
  assign n24504 = ~n6739 & n24503;
  assign n24505 = ~n7945 & n24504;
  assign n24506 = ~n7944 & n24505;
  assign n24507 = ~n7807 & n24506;
  assign n24508 = ~n7943 & n24507;
  assign n24509 = n7966 & n24508;
  assign n24510 = n7942 & n24509;
  assign n24511 = n7935 & n24510;
  assign n24512 = n8264 & n22939;
  assign n24513 = ~n6784 & n24512;
  assign n24514 = ~n8232 & n24513;
  assign n24515 = ~n8017 & n24514;
  assign n24516 = ~n7158 & n24515;
  assign n24517 = ~n8231 & n24516;
  assign n24518 = n8247 & n24517;
  assign n24519 = n8230 & n24518;
  assign n24520 = n8227 & n24519;
  assign n24521 = ~n24511 & ~n24520;
  assign n24522 = n24490 & n24521;
  assign n24523 = n24445 & n24522;
  assign n24524 = ~n1958 & n19228;
  assign n24525 = n7910 & n24524;
  assign n24526 = ~n2242 & n24525;
  assign n24527 = ~n3095 & n24526;
  assign n24528 = ~n3997 & n24527;
  assign n24529 = ~n4003 & n24528;
  assign n24530 = ~n4837 & n24529;
  assign n24531 = ~n5822 & n24530;
  assign n24532 = ~n6820 & n24531;
  assign n24533 = ~n7907 & n24532;
  assign n24534 = ~n7906 & n24533;
  assign n24535 = ~n7785 & n24534;
  assign n24536 = ~n7905 & n24535;
  assign n24537 = n7925 & n24536;
  assign n24538 = n7904 & n24537;
  assign n24539 = n7897 & n24538;
  assign n24540 = n7978 & n22949;
  assign n24541 = ~n3066 & n24540;
  assign n24542 = ~n3983 & n24541;
  assign n24543 = ~n4003 & n24542;
  assign n24544 = ~n4024 & n24543;
  assign n24545 = ~n4999 & n24544;
  assign n24546 = ~n5827 & n24545;
  assign n24547 = ~n7870 & n24546;
  assign n24548 = ~n7842 & n24547;
  assign n24549 = ~n6893 & n24548;
  assign n24550 = ~n7841 & n24549;
  assign n24551 = n7887 & n24550;
  assign n24552 = n7840 & n24551;
  assign n24553 = n7810 & n24552;
  assign n24554 = pi150 & ~n6754;
  assign n24555 = ~n8017 & n24554;
  assign n24556 = ~n7204 & n24555;
  assign n24557 = ~n8282 & n24556;
  assign n24558 = n8288 & n24557;
  assign n24559 = n8281 & n24558;
  assign n24560 = n8280 & n24559;
  assign n24561 = ~n24553 & ~n24560;
  assign n24562 = ~n24539 & n24561;
  assign n24563 = n8121 & n22925;
  assign n24564 = ~n4817 & n24563;
  assign n24565 = ~n4902 & n24564;
  assign n24566 = ~n6001 & n24565;
  assign n24567 = ~n8094 & n24566;
  assign n24568 = ~n8017 & n24567;
  assign n24569 = ~n7014 & n24568;
  assign n24570 = ~n8093 & n24569;
  assign n24571 = n8111 & n24570;
  assign n24572 = n8092 & n24571;
  assign n24573 = n8086 & n24572;
  assign n24574 = pi166 & ~n8391;
  assign n24575 = ~po161 & n24574;
  assign n24576 = ~n8017 & n24575;
  assign n24577 = ~n8314 & n24576;
  assign n24578 = n8281 & n24577;
  assign n24579 = n8390 & n24578;
  assign n24580 = n8383 & n24579;
  assign n24581 = ~n24573 & ~n24580;
  assign n24582 = n8193 & n22899;
  assign n24583 = ~n5808 & n24582;
  assign n24584 = ~n6056 & n24583;
  assign n24585 = ~n8161 & n24584;
  assign n24586 = ~n8017 & n24585;
  assign n24587 = ~n7073 & n24586;
  assign n24588 = ~n8160 & n24587;
  assign n24589 = n8176 & n24588;
  assign n24590 = n8159 & n24589;
  assign n24591 = n8154 & n24590;
  assign n24592 = pi158 & ~n7663;
  assign n24593 = n8360 & n24592;
  assign n24594 = n8368 & n24593;
  assign n24595 = ~n7869 & n24594;
  assign n24596 = ~n8017 & n24595;
  assign n24597 = ~n8045 & n24596;
  assign n24598 = ~n8335 & n24597;
  assign n24599 = n8331 & n24598;
  assign n24600 = n8328 & n24599;
  assign n24601 = n8306 & n24600;
  assign n24602 = ~n24591 & ~n24601;
  assign n24603 = n24581 & n24602;
  assign n24604 = n24562 & n24603;
  assign po095 = ~n24523 | ~n24604;
  assign n24606 = pi167 & ~n8758;
  assign n24607 = ~n8759 & n24606;
  assign n24608 = ~n8757 & n24607;
  assign n24609 = ~n8792 & n24608;
  assign n24610 = n9938 & n24609;
  assign n24611 = n9936 & n24610;
  assign n24612 = n9943 & n24611;
  assign n24613 = ~n8834 & n24612;
  assign n24614 = ~n9185 & n24613;
  assign n24615 = ~n9207 & n24614;
  assign n24616 = ~n9458 & n24615;
  assign n24617 = n9955 & n24616;
  assign n24618 = n9933 & n24617;
  assign n24619 = n10001 & n24618;
  assign n24620 = ~n1208 & n23206;
  assign n24621 = n4920 & n24620;
  assign n24622 = ~n1270 & n24621;
  assign n24623 = n4932 & n24622;
  assign n24624 = ~n1372 & n24623;
  assign n24625 = ~n2243 & n24624;
  assign n24626 = ~n3104 & n24625;
  assign n24627 = ~n3971 & n24626;
  assign n24628 = ~n4003 & n24627;
  assign n24629 = ~n4872 & n24628;
  assign n24630 = ~n5801 & n24629;
  assign n24631 = ~n6739 & n24630;
  assign n24632 = ~n7807 & n24631;
  assign n24633 = ~n9070 & n24632;
  assign n24634 = ~n9069 & n24633;
  assign n24635 = ~n9068 & n24634;
  assign n24636 = ~n9067 & n24635;
  assign n24637 = n9066 & n24636;
  assign n24638 = n9060 & n24637;
  assign n24639 = n9053 & n24638;
  assign n24640 = ~n24619 & ~n24639;
  assign n24641 = ~n5170 & n10602;
  assign n24642 = n23193 & n24641;
  assign n24643 = ~n5808 & n24642;
  assign n24644 = ~n6056 & n24643;
  assign n24645 = ~n7073 & n24644;
  assign n24646 = ~n9330 & n24645;
  assign n24647 = ~n9185 & n24646;
  assign n24648 = ~n8179 & n24647;
  assign n24649 = ~n9329 & n24648;
  assign n24650 = n9328 & n24649;
  assign n24651 = n9323 & n24650;
  assign n24652 = n9316 & n24651;
  assign n24653 = ~n7204 & n23161;
  assign n24654 = ~n9185 & n24653;
  assign n24655 = ~n8291 & n24654;
  assign n24656 = ~n9444 & n24655;
  assign n24657 = n9450 & n24656;
  assign n24658 = n9443 & n24657;
  assign n24659 = n9442 & n24658;
  assign n24660 = ~n24652 & ~n24659;
  assign n24661 = n24640 & n24660;
  assign n24662 = ~n8218 & n23092;
  assign n24663 = ~n9185 & n24662;
  assign n24664 = n9324 & n24663;
  assign n24665 = n9379 & n24664;
  assign n24666 = n9373 & n24665;
  assign n24667 = pi183 & ~n501;
  assign n24668 = n10133 & n24667;
  assign n24669 = n10138 & n24668;
  assign n24670 = n10131 & n24669;
  assign n24671 = ~n1172 & n24670;
  assign n24672 = ~n1114 & n24671;
  assign n24673 = ~n996 & n24672;
  assign n24674 = ~n500 & n24673;
  assign n24675 = n2316 & n24674;
  assign n24676 = n7608 & n24675;
  assign n24677 = n9915 & n24676;
  assign n24678 = n9856 & n24677;
  assign n24679 = n9733 & n24678;
  assign n24680 = ~n7236 & n24679;
  assign n24681 = ~n6137 & n24680;
  assign n24682 = n6193 & n24681;
  assign n24683 = n6134 & n24682;
  assign n24684 = ~n8867 & n24683;
  assign n24685 = ~n7235 & n24684;
  assign n24686 = n7296 & n24685;
  assign n24687 = n7231 & n24686;
  assign n24688 = ~n8866 & n24687;
  assign n24689 = n8898 & n24688;
  assign n24690 = n8863 & n24689;
  assign n24691 = ~n7999 & n23097;
  assign n24692 = ~n9154 & n24691;
  assign n24693 = n9159 & n24692;
  assign n24694 = ~n24690 & ~n24693;
  assign n24695 = ~n24666 & n24694;
  assign n24696 = ~n8145 & n23067;
  assign n24697 = ~n9185 & n24696;
  assign n24698 = ~n9207 & n24697;
  assign n24699 = n9305 & n24698;
  assign n24700 = n9299 & n24699;
  assign n24701 = ~n8053 & n23041;
  assign n24702 = ~n9185 & n24701;
  assign n24703 = ~n9206 & n24702;
  assign n24704 = n9214 & n24703;
  assign n24705 = ~n24700 & ~n24704;
  assign n24706 = n24695 & n24705;
  assign n24707 = pi175 & ~n9511;
  assign n24708 = ~n8900 & n24707;
  assign n24709 = ~n9185 & n24708;
  assign n24710 = ~n9458 & n24709;
  assign n24711 = n9517 & n24710;
  assign n24712 = n9443 & n24711;
  assign n24713 = n9532 & n24712;
  assign n24714 = pi159 & ~po161;
  assign n24715 = ~n9185 & n24714;
  assign n24716 = ~n8397 & n24715;
  assign n24717 = ~n9458 & n24716;
  assign n24718 = n9443 & n24717;
  assign n24719 = n10088 & n24718;
  assign n24720 = n10081 & n24719;
  assign n24721 = ~n24713 & ~n24720;
  assign n24722 = n24706 & n24721;
  assign n24723 = n24661 & n24722;
  assign n24724 = ~n3373 & n11814;
  assign n24725 = ~n3464 & n24724;
  assign n24726 = n23075 & n24725;
  assign n24727 = ~n3940 & n24726;
  assign n24728 = ~n4001 & n24727;
  assign n24729 = ~n5043 & n24728;
  assign n24730 = ~n5943 & n24729;
  assign n24731 = ~n6951 & n24730;
  assign n24732 = ~n9186 & n24731;
  assign n24733 = ~n9185 & n24732;
  assign n24734 = ~n8037 & n24733;
  assign n24735 = ~n9184 & n24734;
  assign n24736 = n9183 & n24735;
  assign n24737 = n9176 & n24736;
  assign n24738 = n9169 & n24737;
  assign n24739 = pi151 & ~n7411;
  assign n24740 = ~n7412 & n24739;
  assign n24741 = ~n7410 & n24740;
  assign n24742 = ~n7663 & n24741;
  assign n24743 = n8358 & n24742;
  assign n24744 = n9496 & n24743;
  assign n24745 = n7357 & ~n7386;
  assign n24746 = ~n7595 & n24745;
  assign n24747 = n24744 & n24746;
  assign n24748 = ~n7869 & n24747;
  assign n24749 = ~n9472 & n24748;
  assign n24750 = ~n9185 & n24749;
  assign n24751 = ~n8346 & n24750;
  assign n24752 = ~n9471 & n24751;
  assign n24753 = n9470 & n24752;
  assign n24754 = n9467 & n24753;
  assign n24755 = n9460 & n24754;
  assign n24756 = n5775 & n23168;
  assign n24757 = ~n3024 & n13319;
  assign n24758 = n24756 & n24757;
  assign n24759 = ~n3066 & n24758;
  assign n24760 = ~n3983 & n24759;
  assign n24761 = ~n4003 & n24760;
  assign n24762 = ~n4024 & n24761;
  assign n24763 = ~n4999 & n24762;
  assign n24764 = ~n5827 & n24763;
  assign n24765 = ~n6893 & n24764;
  assign n24766 = ~n9114 & n24765;
  assign n24767 = ~n9113 & n24766;
  assign n24768 = ~n7890 & n24767;
  assign n24769 = ~n9112 & n24768;
  assign n24770 = n9111 & n24769;
  assign n24771 = n9104 & n24770;
  assign n24772 = n9097 & n24771;
  assign n24773 = ~n24755 & ~n24772;
  assign n24774 = ~n24738 & n24773;
  assign n24775 = ~n1897 & n18466;
  assign n24776 = n1743 & n24775;
  assign n24777 = ~n2242 & n24776;
  assign n24778 = ~n3095 & n24777;
  assign n24779 = ~n3997 & n24778;
  assign n24780 = ~n4003 & n24779;
  assign n24781 = ~n4837 & n24780;
  assign n24782 = ~n5822 & n24781;
  assign n24783 = ~n6820 & n24782;
  assign n24784 = ~n7785 & n24783;
  assign n24785 = ~n9029 & n24784;
  assign n24786 = ~n9028 & n24785;
  assign n24787 = ~n9027 & n24786;
  assign n24788 = ~n9010 & n24787;
  assign n24789 = n9009 & n24788;
  assign n24790 = n9002 & n24789;
  assign n24791 = n8995 & n24790;
  assign n24792 = pi135 & ~n6461;
  assign n24793 = n6343 & n24792;
  assign n24794 = n8233 & n24793;
  assign n24795 = n9425 & n24794;
  assign n24796 = ~n6784 & n24795;
  assign n24797 = ~n7158 & n24796;
  assign n24798 = ~n9402 & n24797;
  assign n24799 = ~n9185 & n24798;
  assign n24800 = ~n8250 & n24799;
  assign n24801 = ~n9401 & n24800;
  assign n24802 = n9400 & n24801;
  assign n24803 = n9397 & n24802;
  assign n24804 = n9390 & n24803;
  assign n24805 = ~n24791 & ~n24804;
  assign n24806 = n9282 & n20698;
  assign n24807 = ~n4817 & n24806;
  assign n24808 = ~n4902 & n24807;
  assign n24809 = ~n6001 & n24808;
  assign n24810 = ~n7014 & n24809;
  assign n24811 = ~n9261 & n24810;
  assign n24812 = ~n9185 & n24811;
  assign n24813 = ~n8114 & n24812;
  assign n24814 = ~n9260 & n24813;
  assign n24815 = n9259 & n24814;
  assign n24816 = n9253 & n24815;
  assign n24817 = n9246 & n24816;
  assign n24818 = pi191 & ~n501;
  assign n24819 = n5714 & n24818;
  assign n24820 = n5719 & n24819;
  assign n24821 = n8912 & n24820;
  assign n24822 = ~n1172 & n24821;
  assign n24823 = ~n996 & n24822;
  assign n24824 = ~n2306 & n24823;
  assign n24825 = ~n500 & n24824;
  assign n24826 = n2316 & n24825;
  assign n24827 = n7608 & n24826;
  assign n24828 = n10030 & n24827;
  assign n24829 = n10029 & n24828;
  assign n24830 = ~n7236 & n24829;
  assign n24831 = ~n6137 & n24830;
  assign n24832 = n6193 & n24831;
  assign n24833 = n6134 & n24832;
  assign n24834 = ~n8867 & n24833;
  assign n24835 = ~n7235 & n24834;
  assign n24836 = n7296 & n24835;
  assign n24837 = n7231 & n24836;
  assign n24838 = ~n10027 & n24837;
  assign n24839 = ~n8866 & n24838;
  assign n24840 = n8898 & n24839;
  assign n24841 = n8863 & n24840;
  assign n24842 = ~n10026 & n24841;
  assign n24843 = n10072 & n24842;
  assign n24844 = n10021 & n24843;
  assign n24845 = ~n24817 & ~n24844;
  assign n24846 = n24805 & n24845;
  assign n24847 = n24774 & n24846;
  assign po096 = ~n24723 | ~n24847;
  assign n24849 = n8358 & n23403;
  assign n24850 = n9496 & n24849;
  assign n24851 = n9499 & n24850;
  assign n24852 = ~n7869 & n24851;
  assign n24853 = ~n9472 & n24852;
  assign n24854 = ~n9185 & n24853;
  assign n24855 = ~n8346 & n24854;
  assign n24856 = ~n9471 & n24855;
  assign n24857 = n9470 & n24856;
  assign n24858 = n9467 & n24857;
  assign n24859 = n9460 & n24858;
  assign n24860 = n3846 & n21883;
  assign n24861 = n3854 & n24860;
  assign n24862 = n9138 & n24861;
  assign n24863 = ~n3066 & n24862;
  assign n24864 = ~n3983 & n24863;
  assign n24865 = ~n4003 & n24864;
  assign n24866 = ~n4024 & n24865;
  assign n24867 = ~n4999 & n24866;
  assign n24868 = ~n5827 & n24867;
  assign n24869 = ~n6893 & n24868;
  assign n24870 = ~n9114 & n24869;
  assign n24871 = ~n9113 & n24870;
  assign n24872 = ~n7890 & n24871;
  assign n24873 = ~n9112 & n24872;
  assign n24874 = n9111 & n24873;
  assign n24875 = n9104 & n24874;
  assign n24876 = n9097 & n24875;
  assign n24877 = ~n24859 & ~n24876;
  assign n24878 = pi136 & ~n6461;
  assign n24879 = n6343 & n24878;
  assign n24880 = n8233 & n24879;
  assign n24881 = n9425 & n24880;
  assign n24882 = ~n6784 & n24881;
  assign n24883 = ~n7158 & n24882;
  assign n24884 = ~n9402 & n24883;
  assign n24885 = ~n9185 & n24884;
  assign n24886 = ~n8250 & n24885;
  assign n24887 = ~n9401 & n24886;
  assign n24888 = n9400 & n24887;
  assign n24889 = n9397 & n24888;
  assign n24890 = n9390 & n24889;
  assign n24891 = ~n1208 & n23366;
  assign n24892 = n4920 & n24891;
  assign n24893 = ~n1270 & n24892;
  assign n24894 = n4932 & n24893;
  assign n24895 = ~n1372 & n24894;
  assign n24896 = ~n2243 & n24895;
  assign n24897 = ~n3104 & n24896;
  assign n24898 = ~n3971 & n24897;
  assign n24899 = ~n4003 & n24898;
  assign n24900 = ~n4872 & n24899;
  assign n24901 = ~n5801 & n24900;
  assign n24902 = ~n6739 & n24901;
  assign n24903 = ~n7807 & n24902;
  assign n24904 = ~n9070 & n24903;
  assign n24905 = ~n9069 & n24904;
  assign n24906 = ~n9068 & n24905;
  assign n24907 = ~n9067 & n24906;
  assign n24908 = n9066 & n24907;
  assign n24909 = n9060 & n24908;
  assign n24910 = n9053 & n24909;
  assign n24911 = ~n24890 & ~n24910;
  assign n24912 = n24877 & n24911;
  assign n24913 = ~n8053 & n23255;
  assign n24914 = ~n9185 & n24913;
  assign n24915 = ~n9206 & n24914;
  assign n24916 = n9214 & n24915;
  assign n24917 = pi184 & ~n501;
  assign n24918 = n10133 & n24917;
  assign n24919 = n10138 & n24918;
  assign n24920 = n10131 & n24919;
  assign n24921 = ~n1172 & n24920;
  assign n24922 = ~n1114 & n24921;
  assign n24923 = ~n996 & n24922;
  assign n24924 = ~n500 & n24923;
  assign n24925 = n2316 & n24924;
  assign n24926 = n7608 & n24925;
  assign n24927 = n9915 & n24926;
  assign n24928 = n9856 & n24927;
  assign n24929 = n9733 & n24928;
  assign n24930 = ~n7236 & n24929;
  assign n24931 = ~n6137 & n24930;
  assign n24932 = n6193 & n24931;
  assign n24933 = n6134 & n24932;
  assign n24934 = ~n8867 & n24933;
  assign n24935 = ~n7235 & n24934;
  assign n24936 = n7296 & n24935;
  assign n24937 = n7231 & n24936;
  assign n24938 = ~n8866 & n24937;
  assign n24939 = n8898 & n24938;
  assign n24940 = n8863 & n24939;
  assign n24941 = ~n7999 & n23304;
  assign n24942 = ~n9154 & n24941;
  assign n24943 = n9159 & n24942;
  assign n24944 = ~n24940 & ~n24943;
  assign n24945 = ~n24916 & n24944;
  assign n24946 = ~n8145 & n23299;
  assign n24947 = ~n9185 & n24946;
  assign n24948 = ~n9207 & n24947;
  assign n24949 = n9305 & n24948;
  assign n24950 = n9299 & n24949;
  assign n24951 = ~n8218 & n23260;
  assign n24952 = ~n9185 & n24951;
  assign n24953 = n9324 & n24952;
  assign n24954 = n9379 & n24953;
  assign n24955 = n9373 & n24954;
  assign n24956 = ~n24950 & ~n24955;
  assign n24957 = n24945 & n24956;
  assign n24958 = n9282 & n20846;
  assign n24959 = ~n4817 & n24958;
  assign n24960 = ~n4902 & n24959;
  assign n24961 = ~n6001 & n24960;
  assign n24962 = ~n7014 & n24961;
  assign n24963 = ~n9261 & n24962;
  assign n24964 = ~n9185 & n24963;
  assign n24965 = ~n8114 & n24964;
  assign n24966 = ~n9260 & n24965;
  assign n24967 = n9259 & n24966;
  assign n24968 = n9253 & n24967;
  assign n24969 = n9246 & n24968;
  assign n24970 = pi168 & ~n8762;
  assign n24971 = n8822 & n24970;
  assign n24972 = n8664 & n24971;
  assign n24973 = n10172 & n24972;
  assign n24974 = ~n8834 & n24973;
  assign n24975 = ~n9185 & n24974;
  assign n24976 = ~n9207 & n24975;
  assign n24977 = ~n9458 & n24976;
  assign n24978 = n9955 & n24977;
  assign n24979 = n9933 & n24978;
  assign n24980 = n10001 & n24979;
  assign n24981 = ~n24969 & ~n24980;
  assign n24982 = n24957 & n24981;
  assign n24983 = n24912 & n24982;
  assign n24984 = n3740 & n19386;
  assign n24985 = n3951 & n24984;
  assign n24986 = n9220 & n24985;
  assign n24987 = ~n3940 & n24986;
  assign n24988 = ~n4001 & n24987;
  assign n24989 = ~n5043 & n24988;
  assign n24990 = ~n5943 & n24989;
  assign n24991 = ~n6951 & n24990;
  assign n24992 = ~n9186 & n24991;
  assign n24993 = ~n9185 & n24992;
  assign n24994 = ~n8037 & n24993;
  assign n24995 = ~n9184 & n24994;
  assign n24996 = n9183 & n24995;
  assign n24997 = n9176 & n24996;
  assign n24998 = n9169 & n24997;
  assign n24999 = pi160 & ~po161;
  assign n25000 = ~n9185 & n24999;
  assign n25001 = ~n8397 & n25000;
  assign n25002 = ~n9458 & n25001;
  assign n25003 = n9443 & n25002;
  assign n25004 = n10088 & n25003;
  assign n25005 = n10081 & n25004;
  assign n25006 = pi176 & ~n9511;
  assign n25007 = ~n8900 & n25006;
  assign n25008 = ~n9185 & n25007;
  assign n25009 = ~n9458 & n25008;
  assign n25010 = n9517 & n25009;
  assign n25011 = n9443 & n25010;
  assign n25012 = n9532 & n25011;
  assign n25013 = ~n25005 & ~n25012;
  assign n25014 = ~n24998 & n25013;
  assign n25015 = ~n1897 & n18504;
  assign n25016 = n1743 & n25015;
  assign n25017 = ~n2242 & n25016;
  assign n25018 = ~n3095 & n25017;
  assign n25019 = ~n3997 & n25018;
  assign n25020 = ~n4003 & n25019;
  assign n25021 = ~n4837 & n25020;
  assign n25022 = ~n5822 & n25021;
  assign n25023 = ~n6820 & n25022;
  assign n25024 = ~n7785 & n25023;
  assign n25025 = ~n9029 & n25024;
  assign n25026 = ~n9028 & n25025;
  assign n25027 = ~n9027 & n25026;
  assign n25028 = ~n9010 & n25027;
  assign n25029 = n9009 & n25028;
  assign n25030 = n9002 & n25029;
  assign n25031 = n8995 & n25030;
  assign n25032 = pi192 & ~n501;
  assign n25033 = n5714 & n25032;
  assign n25034 = n5719 & n25033;
  assign n25035 = n8912 & n25034;
  assign n25036 = ~n1172 & n25035;
  assign n25037 = ~n996 & n25036;
  assign n25038 = ~n2306 & n25037;
  assign n25039 = ~n500 & n25038;
  assign n25040 = n2316 & n25039;
  assign n25041 = n7608 & n25040;
  assign n25042 = n10030 & n25041;
  assign n25043 = n10029 & n25042;
  assign n25044 = ~n7236 & n25043;
  assign n25045 = ~n6137 & n25044;
  assign n25046 = n6193 & n25045;
  assign n25047 = n6134 & n25046;
  assign n25048 = ~n8867 & n25047;
  assign n25049 = ~n7235 & n25048;
  assign n25050 = n7296 & n25049;
  assign n25051 = n7231 & n25050;
  assign n25052 = ~n10027 & n25051;
  assign n25053 = ~n8866 & n25052;
  assign n25054 = n8898 & n25053;
  assign n25055 = n8863 & n25054;
  assign n25056 = ~n10026 & n25055;
  assign n25057 = n10072 & n25056;
  assign n25058 = n10021 & n25057;
  assign n25059 = ~n25031 & ~n25058;
  assign n25060 = ~n7204 & n23413;
  assign n25061 = ~n9185 & n25060;
  assign n25062 = ~n8291 & n25061;
  assign n25063 = ~n9444 & n25062;
  assign n25064 = n9450 & n25063;
  assign n25065 = n9443 & n25064;
  assign n25066 = n9442 & n25065;
  assign n25067 = n9355 & n20901;
  assign n25068 = ~n5808 & n25067;
  assign n25069 = ~n6056 & n25068;
  assign n25070 = ~n7073 & n25069;
  assign n25071 = ~n9330 & n25070;
  assign n25072 = ~n9185 & n25071;
  assign n25073 = ~n8179 & n25072;
  assign n25074 = ~n9329 & n25073;
  assign n25075 = n9328 & n25074;
  assign n25076 = n9323 & n25075;
  assign n25077 = n9316 & n25076;
  assign n25078 = ~n25066 & ~n25077;
  assign n25079 = n25059 & n25078;
  assign n25080 = n25014 & n25079;
  assign po097 = ~n24983 | ~n25080;
  assign n25082 = ~n1897 & n18542;
  assign n25083 = n1743 & n25082;
  assign n25084 = ~n2242 & n25083;
  assign n25085 = ~n3095 & n25084;
  assign n25086 = ~n3997 & n25085;
  assign n25087 = ~n4003 & n25086;
  assign n25088 = ~n4837 & n25087;
  assign n25089 = ~n5822 & n25088;
  assign n25090 = ~n6820 & n25089;
  assign n25091 = ~n7785 & n25090;
  assign n25092 = ~n9029 & n25091;
  assign n25093 = ~n9028 & n25092;
  assign n25094 = ~n9027 & n25093;
  assign n25095 = ~n9010 & n25094;
  assign n25096 = n9009 & n25095;
  assign n25097 = n9002 & n25096;
  assign n25098 = n8995 & n25097;
  assign n25099 = pi193 & ~n501;
  assign n25100 = n5714 & n25099;
  assign n25101 = n5719 & n25100;
  assign n25102 = n8912 & n25101;
  assign n25103 = ~n1172 & n25102;
  assign n25104 = ~n996 & n25103;
  assign n25105 = ~n2306 & n25104;
  assign n25106 = ~n500 & n25105;
  assign n25107 = n2316 & n25106;
  assign n25108 = n7608 & n25107;
  assign n25109 = n10030 & n25108;
  assign n25110 = n10029 & n25109;
  assign n25111 = ~n7236 & n25110;
  assign n25112 = ~n6137 & n25111;
  assign n25113 = n6193 & n25112;
  assign n25114 = n6134 & n25113;
  assign n25115 = ~n8867 & n25114;
  assign n25116 = ~n7235 & n25115;
  assign n25117 = n7296 & n25116;
  assign n25118 = n7231 & n25117;
  assign n25119 = ~n10027 & n25118;
  assign n25120 = ~n8866 & n25119;
  assign n25121 = n8898 & n25120;
  assign n25122 = n8863 & n25121;
  assign n25123 = ~n10026 & n25122;
  assign n25124 = n10072 & n25123;
  assign n25125 = n10021 & n25124;
  assign n25126 = ~n25098 & ~n25125;
  assign n25127 = pi161 & ~po161;
  assign n25128 = ~n9185 & n25127;
  assign n25129 = ~n8397 & n25128;
  assign n25130 = ~n9458 & n25129;
  assign n25131 = n9443 & n25130;
  assign n25132 = n10088 & n25131;
  assign n25133 = n10081 & n25132;
  assign n25134 = pi137 & ~n6461;
  assign n25135 = n6343 & n25134;
  assign n25136 = n8233 & n25135;
  assign n25137 = n9425 & n25136;
  assign n25138 = ~n6784 & n25137;
  assign n25139 = ~n7158 & n25138;
  assign n25140 = ~n9402 & n25139;
  assign n25141 = ~n9185 & n25140;
  assign n25142 = ~n8250 & n25141;
  assign n25143 = ~n9401 & n25142;
  assign n25144 = n9400 & n25143;
  assign n25145 = n9397 & n25144;
  assign n25146 = n9390 & n25145;
  assign n25147 = ~n25133 & ~n25146;
  assign n25148 = n25126 & n25147;
  assign n25149 = ~n8145 & n23470;
  assign n25150 = ~n9185 & n25149;
  assign n25151 = ~n9207 & n25150;
  assign n25152 = n9305 & n25151;
  assign n25153 = n9299 & n25152;
  assign n25154 = ~n7999 & n23499;
  assign n25155 = ~n9154 & n25154;
  assign n25156 = n9159 & n25155;
  assign n25157 = pi185 & ~n501;
  assign n25158 = n10133 & n25157;
  assign n25159 = n10138 & n25158;
  assign n25160 = n10131 & n25159;
  assign n25161 = ~n1172 & n25160;
  assign n25162 = ~n1114 & n25161;
  assign n25163 = ~n996 & n25162;
  assign n25164 = ~n500 & n25163;
  assign n25165 = n2316 & n25164;
  assign n25166 = n7608 & n25165;
  assign n25167 = n9915 & n25166;
  assign n25168 = n9856 & n25167;
  assign n25169 = n9733 & n25168;
  assign n25170 = ~n7236 & n25169;
  assign n25171 = ~n6137 & n25170;
  assign n25172 = n6193 & n25171;
  assign n25173 = n6134 & n25172;
  assign n25174 = ~n8867 & n25173;
  assign n25175 = ~n7235 & n25174;
  assign n25176 = n7296 & n25175;
  assign n25177 = n7231 & n25176;
  assign n25178 = ~n8866 & n25177;
  assign n25179 = n8898 & n25178;
  assign n25180 = n8863 & n25179;
  assign n25181 = ~n25156 & ~n25180;
  assign n25182 = ~n25153 & n25181;
  assign n25183 = ~n8053 & n23495;
  assign n25184 = ~n9185 & n25183;
  assign n25185 = ~n9206 & n25184;
  assign n25186 = n9214 & n25185;
  assign n25187 = ~n8218 & n23476;
  assign n25188 = ~n9185 & n25187;
  assign n25189 = n9324 & n25188;
  assign n25190 = n9379 & n25189;
  assign n25191 = n9373 & n25190;
  assign n25192 = ~n25186 & ~n25191;
  assign n25193 = n25182 & n25192;
  assign n25194 = n9282 & n21037;
  assign n25195 = ~n4817 & n25194;
  assign n25196 = ~n4902 & n25195;
  assign n25197 = ~n6001 & n25196;
  assign n25198 = ~n7014 & n25197;
  assign n25199 = ~n9261 & n25198;
  assign n25200 = ~n9185 & n25199;
  assign n25201 = ~n8114 & n25200;
  assign n25202 = ~n9260 & n25201;
  assign n25203 = n9259 & n25202;
  assign n25204 = n9253 & n25203;
  assign n25205 = n9246 & n25204;
  assign n25206 = n3846 & n22055;
  assign n25207 = n3854 & n25206;
  assign n25208 = n9138 & n25207;
  assign n25209 = ~n3066 & n25208;
  assign n25210 = ~n3983 & n25209;
  assign n25211 = ~n4003 & n25210;
  assign n25212 = ~n4024 & n25211;
  assign n25213 = ~n4999 & n25212;
  assign n25214 = ~n5827 & n25213;
  assign n25215 = ~n6893 & n25214;
  assign n25216 = ~n9114 & n25215;
  assign n25217 = ~n9113 & n25216;
  assign n25218 = ~n7890 & n25217;
  assign n25219 = ~n9112 & n25218;
  assign n25220 = n9111 & n25219;
  assign n25221 = n9104 & n25220;
  assign n25222 = n9097 & n25221;
  assign n25223 = ~n25205 & ~n25222;
  assign n25224 = n25193 & n25223;
  assign n25225 = n25148 & n25224;
  assign n25226 = n8358 & n23526;
  assign n25227 = n9496 & n25226;
  assign n25228 = n9499 & n25227;
  assign n25229 = ~n7869 & n25228;
  assign n25230 = ~n9472 & n25229;
  assign n25231 = ~n9185 & n25230;
  assign n25232 = ~n8346 & n25231;
  assign n25233 = ~n9471 & n25232;
  assign n25234 = n9470 & n25233;
  assign n25235 = n9467 & n25234;
  assign n25236 = n9460 & n25235;
  assign n25237 = pi177 & ~n9511;
  assign n25238 = ~n8900 & n25237;
  assign n25239 = ~n9185 & n25238;
  assign n25240 = ~n9458 & n25239;
  assign n25241 = n9517 & n25240;
  assign n25242 = n9443 & n25241;
  assign n25243 = n9532 & n25242;
  assign n25244 = ~n7204 & n23565;
  assign n25245 = ~n9185 & n25244;
  assign n25246 = ~n8291 & n25245;
  assign n25247 = ~n9444 & n25246;
  assign n25248 = n9450 & n25247;
  assign n25249 = n9443 & n25248;
  assign n25250 = n9442 & n25249;
  assign n25251 = ~n25243 & ~n25250;
  assign n25252 = ~n25236 & n25251;
  assign n25253 = pi169 & ~n8762;
  assign n25254 = n8822 & n25253;
  assign n25255 = n8664 & n25254;
  assign n25256 = n10172 & n25255;
  assign n25257 = ~n8834 & n25256;
  assign n25258 = ~n9185 & n25257;
  assign n25259 = ~n9207 & n25258;
  assign n25260 = ~n9458 & n25259;
  assign n25261 = n9955 & n25260;
  assign n25262 = n9933 & n25261;
  assign n25263 = n10001 & n25262;
  assign n25264 = n3740 & n19437;
  assign n25265 = n3951 & n25264;
  assign n25266 = n9220 & n25265;
  assign n25267 = ~n3940 & n25266;
  assign n25268 = ~n4001 & n25267;
  assign n25269 = ~n5043 & n25268;
  assign n25270 = ~n5943 & n25269;
  assign n25271 = ~n6951 & n25270;
  assign n25272 = ~n9186 & n25271;
  assign n25273 = ~n9185 & n25272;
  assign n25274 = ~n8037 & n25273;
  assign n25275 = ~n9184 & n25274;
  assign n25276 = n9183 & n25275;
  assign n25277 = n9176 & n25276;
  assign n25278 = n9169 & n25277;
  assign n25279 = ~n25263 & ~n25278;
  assign n25280 = ~n1208 & n23616;
  assign n25281 = n4920 & n25280;
  assign n25282 = ~n1270 & n25281;
  assign n25283 = n4932 & n25282;
  assign n25284 = ~n1372 & n25283;
  assign n25285 = ~n2243 & n25284;
  assign n25286 = ~n3104 & n25285;
  assign n25287 = ~n3971 & n25286;
  assign n25288 = ~n4003 & n25287;
  assign n25289 = ~n4872 & n25288;
  assign n25290 = ~n5801 & n25289;
  assign n25291 = ~n6739 & n25290;
  assign n25292 = ~n7807 & n25291;
  assign n25293 = ~n9070 & n25292;
  assign n25294 = ~n9069 & n25293;
  assign n25295 = ~n9068 & n25294;
  assign n25296 = ~n9067 & n25295;
  assign n25297 = n9066 & n25296;
  assign n25298 = n9060 & n25297;
  assign n25299 = n9053 & n25298;
  assign n25300 = n9355 & n21027;
  assign n25301 = ~n5808 & n25300;
  assign n25302 = ~n6056 & n25301;
  assign n25303 = ~n7073 & n25302;
  assign n25304 = ~n9330 & n25303;
  assign n25305 = ~n9185 & n25304;
  assign n25306 = ~n8179 & n25305;
  assign n25307 = ~n9329 & n25306;
  assign n25308 = n9328 & n25307;
  assign n25309 = n9323 & n25308;
  assign n25310 = n9316 & n25309;
  assign n25311 = ~n25299 & ~n25310;
  assign n25312 = n25279 & n25311;
  assign n25313 = n25252 & n25312;
  assign po098 = ~n25225 | ~n25313;
  assign n25315 = pi162 & ~po161;
  assign n25316 = ~n9185 & n25315;
  assign n25317 = ~n8397 & n25316;
  assign n25318 = ~n9458 & n25317;
  assign n25319 = n9443 & n25318;
  assign n25320 = n10088 & n25319;
  assign n25321 = n10081 & n25320;
  assign n25322 = ~n1897 & n18580;
  assign n25323 = n1743 & n25322;
  assign n25324 = ~n2242 & n25323;
  assign n25325 = ~n3095 & n25324;
  assign n25326 = ~n3997 & n25325;
  assign n25327 = ~n4003 & n25326;
  assign n25328 = ~n4837 & n25327;
  assign n25329 = ~n5822 & n25328;
  assign n25330 = ~n6820 & n25329;
  assign n25331 = ~n7785 & n25330;
  assign n25332 = ~n9029 & n25331;
  assign n25333 = ~n9028 & n25332;
  assign n25334 = ~n9027 & n25333;
  assign n25335 = ~n9010 & n25334;
  assign n25336 = n9009 & n25335;
  assign n25337 = n9002 & n25336;
  assign n25338 = n8995 & n25337;
  assign n25339 = ~n25321 & ~n25338;
  assign n25340 = pi178 & ~n9511;
  assign n25341 = ~n8900 & n25340;
  assign n25342 = ~n9185 & n25341;
  assign n25343 = ~n9458 & n25342;
  assign n25344 = n9517 & n25343;
  assign n25345 = n9443 & n25344;
  assign n25346 = n9532 & n25345;
  assign n25347 = ~n7204 & n23781;
  assign n25348 = ~n9185 & n25347;
  assign n25349 = ~n8291 & n25348;
  assign n25350 = ~n9444 & n25349;
  assign n25351 = n9450 & n25350;
  assign n25352 = n9443 & n25351;
  assign n25353 = n9442 & n25352;
  assign n25354 = ~n25346 & ~n25353;
  assign n25355 = n25339 & n25354;
  assign n25356 = ~n8145 & n23651;
  assign n25357 = ~n9185 & n25356;
  assign n25358 = ~n9207 & n25357;
  assign n25359 = n9305 & n25358;
  assign n25360 = n9299 & n25359;
  assign n25361 = ~n7999 & n23692;
  assign n25362 = ~n9154 & n25361;
  assign n25363 = n9159 & n25362;
  assign n25364 = pi186 & ~n501;
  assign n25365 = n10133 & n25364;
  assign n25366 = n10138 & n25365;
  assign n25367 = n10131 & n25366;
  assign n25368 = ~n1172 & n25367;
  assign n25369 = ~n1114 & n25368;
  assign n25370 = ~n996 & n25369;
  assign n25371 = ~n500 & n25370;
  assign n25372 = n2316 & n25371;
  assign n25373 = n7608 & n25372;
  assign n25374 = n9915 & n25373;
  assign n25375 = n9856 & n25374;
  assign n25376 = n9733 & n25375;
  assign n25377 = ~n7236 & n25376;
  assign n25378 = ~n6137 & n25377;
  assign n25379 = n6193 & n25378;
  assign n25380 = n6134 & n25379;
  assign n25381 = ~n8867 & n25380;
  assign n25382 = ~n7235 & n25381;
  assign n25383 = n7296 & n25382;
  assign n25384 = n7231 & n25383;
  assign n25385 = ~n8866 & n25384;
  assign n25386 = n8898 & n25385;
  assign n25387 = n8863 & n25386;
  assign n25388 = ~n25363 & ~n25387;
  assign n25389 = ~n25360 & n25388;
  assign n25390 = ~n8053 & n23641;
  assign n25391 = ~n9185 & n25390;
  assign n25392 = ~n9206 & n25391;
  assign n25393 = n9214 & n25392;
  assign n25394 = ~n8218 & n23646;
  assign n25395 = ~n9185 & n25394;
  assign n25396 = n9324 & n25395;
  assign n25397 = n9379 & n25396;
  assign n25398 = n9373 & n25397;
  assign n25399 = ~n25393 & ~n25398;
  assign n25400 = n25389 & n25399;
  assign n25401 = n9282 & n21163;
  assign n25402 = ~n4817 & n25401;
  assign n25403 = ~n4902 & n25402;
  assign n25404 = ~n6001 & n25403;
  assign n25405 = ~n7014 & n25404;
  assign n25406 = ~n9261 & n25405;
  assign n25407 = ~n9185 & n25406;
  assign n25408 = ~n8114 & n25407;
  assign n25409 = ~n9260 & n25408;
  assign n25410 = n9259 & n25409;
  assign n25411 = n9253 & n25410;
  assign n25412 = n9246 & n25411;
  assign n25413 = n3846 & n22280;
  assign n25414 = n3854 & n25413;
  assign n25415 = n9138 & n25414;
  assign n25416 = ~n3066 & n25415;
  assign n25417 = ~n3983 & n25416;
  assign n25418 = ~n4003 & n25417;
  assign n25419 = ~n4024 & n25418;
  assign n25420 = ~n4999 & n25419;
  assign n25421 = ~n5827 & n25420;
  assign n25422 = ~n6893 & n25421;
  assign n25423 = ~n9114 & n25422;
  assign n25424 = ~n9113 & n25423;
  assign n25425 = ~n7890 & n25424;
  assign n25426 = ~n9112 & n25425;
  assign n25427 = n9111 & n25426;
  assign n25428 = n9104 & n25427;
  assign n25429 = n9097 & n25428;
  assign n25430 = ~n25412 & ~n25429;
  assign n25431 = n25400 & n25430;
  assign n25432 = n25355 & n25431;
  assign n25433 = pi138 & ~n6461;
  assign n25434 = n6343 & n25433;
  assign n25435 = n8233 & n25434;
  assign n25436 = n9425 & n25435;
  assign n25437 = ~n6784 & n25436;
  assign n25438 = ~n7158 & n25437;
  assign n25439 = ~n9402 & n25438;
  assign n25440 = ~n9185 & n25439;
  assign n25441 = ~n8250 & n25440;
  assign n25442 = ~n9401 & n25441;
  assign n25443 = n9400 & n25442;
  assign n25444 = n9397 & n25443;
  assign n25445 = n9390 & n25444;
  assign n25446 = n9355 & n21153;
  assign n25447 = ~n5808 & n25446;
  assign n25448 = ~n6056 & n25447;
  assign n25449 = ~n7073 & n25448;
  assign n25450 = ~n9330 & n25449;
  assign n25451 = ~n9185 & n25450;
  assign n25452 = ~n8179 & n25451;
  assign n25453 = ~n9329 & n25452;
  assign n25454 = n9328 & n25453;
  assign n25455 = n9323 & n25454;
  assign n25456 = n9316 & n25455;
  assign n25457 = n8358 & n23752;
  assign n25458 = n9496 & n25457;
  assign n25459 = n9499 & n25458;
  assign n25460 = ~n7869 & n25459;
  assign n25461 = ~n9472 & n25460;
  assign n25462 = ~n9185 & n25461;
  assign n25463 = ~n8346 & n25462;
  assign n25464 = ~n9471 & n25463;
  assign n25465 = n9470 & n25464;
  assign n25466 = n9467 & n25465;
  assign n25467 = n9460 & n25466;
  assign n25468 = ~n25456 & ~n25467;
  assign n25469 = ~n25445 & n25468;
  assign n25470 = n3740 & n19508;
  assign n25471 = n3951 & n25470;
  assign n25472 = n9220 & n25471;
  assign n25473 = ~n3940 & n25472;
  assign n25474 = ~n4001 & n25473;
  assign n25475 = ~n5043 & n25474;
  assign n25476 = ~n5943 & n25475;
  assign n25477 = ~n6951 & n25476;
  assign n25478 = ~n9186 & n25477;
  assign n25479 = ~n9185 & n25478;
  assign n25480 = ~n8037 & n25479;
  assign n25481 = ~n9184 & n25480;
  assign n25482 = n9183 & n25481;
  assign n25483 = n9176 & n25482;
  assign n25484 = n9169 & n25483;
  assign n25485 = pi194 & ~n501;
  assign n25486 = n5714 & n25485;
  assign n25487 = n5719 & n25486;
  assign n25488 = n8912 & n25487;
  assign n25489 = ~n1172 & n25488;
  assign n25490 = ~n996 & n25489;
  assign n25491 = ~n2306 & n25490;
  assign n25492 = ~n500 & n25491;
  assign n25493 = n2316 & n25492;
  assign n25494 = n7608 & n25493;
  assign n25495 = n10030 & n25494;
  assign n25496 = n10029 & n25495;
  assign n25497 = ~n7236 & n25496;
  assign n25498 = ~n6137 & n25497;
  assign n25499 = n6193 & n25498;
  assign n25500 = n6134 & n25499;
  assign n25501 = ~n8867 & n25500;
  assign n25502 = ~n7235 & n25501;
  assign n25503 = n7296 & n25502;
  assign n25504 = n7231 & n25503;
  assign n25505 = ~n10027 & n25504;
  assign n25506 = ~n8866 & n25505;
  assign n25507 = n8898 & n25506;
  assign n25508 = n8863 & n25507;
  assign n25509 = ~n10026 & n25508;
  assign n25510 = n10072 & n25509;
  assign n25511 = n10021 & n25510;
  assign n25512 = ~n25484 & ~n25511;
  assign n25513 = pi170 & ~n8762;
  assign n25514 = n8822 & n25513;
  assign n25515 = n8664 & n25514;
  assign n25516 = n10172 & n25515;
  assign n25517 = ~n8834 & n25516;
  assign n25518 = ~n9185 & n25517;
  assign n25519 = ~n9207 & n25518;
  assign n25520 = ~n9458 & n25519;
  assign n25521 = n9955 & n25520;
  assign n25522 = n9933 & n25521;
  assign n25523 = n10001 & n25522;
  assign n25524 = ~n1208 & n23719;
  assign n25525 = n4920 & n25524;
  assign n25526 = ~n1270 & n25525;
  assign n25527 = n4932 & n25526;
  assign n25528 = ~n1372 & n25527;
  assign n25529 = ~n2243 & n25528;
  assign n25530 = ~n3104 & n25529;
  assign n25531 = ~n3971 & n25530;
  assign n25532 = ~n4003 & n25531;
  assign n25533 = ~n4872 & n25532;
  assign n25534 = ~n5801 & n25533;
  assign n25535 = ~n6739 & n25534;
  assign n25536 = ~n7807 & n25535;
  assign n25537 = ~n9070 & n25536;
  assign n25538 = ~n9069 & n25537;
  assign n25539 = ~n9068 & n25538;
  assign n25540 = ~n9067 & n25539;
  assign n25541 = n9066 & n25540;
  assign n25542 = n9060 & n25541;
  assign n25543 = n9053 & n25542;
  assign n25544 = ~n25523 & ~n25543;
  assign n25545 = n25512 & n25544;
  assign n25546 = n25469 & n25545;
  assign po099 = ~n25432 | ~n25546;
  assign n25548 = pi195 & ~n501;
  assign n25549 = n5714 & n25548;
  assign n25550 = n5719 & n25549;
  assign n25551 = n8912 & n25550;
  assign n25552 = ~n1172 & n25551;
  assign n25553 = ~n996 & n25552;
  assign n25554 = ~n2306 & n25553;
  assign n25555 = ~n500 & n25554;
  assign n25556 = n2316 & n25555;
  assign n25557 = n7608 & n25556;
  assign n25558 = n10030 & n25557;
  assign n25559 = n10029 & n25558;
  assign n25560 = ~n7236 & n25559;
  assign n25561 = ~n6137 & n25560;
  assign n25562 = n6193 & n25561;
  assign n25563 = n6134 & n25562;
  assign n25564 = ~n8867 & n25563;
  assign n25565 = ~n7235 & n25564;
  assign n25566 = n7296 & n25565;
  assign n25567 = n7231 & n25566;
  assign n25568 = ~n10027 & n25567;
  assign n25569 = ~n8866 & n25568;
  assign n25570 = n8898 & n25569;
  assign n25571 = n8863 & n25570;
  assign n25572 = ~n10026 & n25571;
  assign n25573 = n10072 & n25572;
  assign n25574 = n10021 & n25573;
  assign n25575 = n8358 & n23945;
  assign n25576 = n9496 & n25575;
  assign n25577 = n9499 & n25576;
  assign n25578 = ~n7869 & n25577;
  assign n25579 = ~n9472 & n25578;
  assign n25580 = ~n9185 & n25579;
  assign n25581 = ~n8346 & n25580;
  assign n25582 = ~n9471 & n25581;
  assign n25583 = n9470 & n25582;
  assign n25584 = n9467 & n25583;
  assign n25585 = n9460 & n25584;
  assign n25586 = ~n25574 & ~n25585;
  assign n25587 = pi139 & ~n6461;
  assign n25588 = n6343 & n25587;
  assign n25589 = n8233 & n25588;
  assign n25590 = n9425 & n25589;
  assign n25591 = ~n6784 & n25590;
  assign n25592 = ~n7158 & n25591;
  assign n25593 = ~n9402 & n25592;
  assign n25594 = ~n9185 & n25593;
  assign n25595 = ~n8250 & n25594;
  assign n25596 = ~n9401 & n25595;
  assign n25597 = n9400 & n25596;
  assign n25598 = n9397 & n25597;
  assign n25599 = n9390 & n25598;
  assign n25600 = pi171 & ~n8762;
  assign n25601 = n8822 & n25600;
  assign n25602 = n8664 & n25601;
  assign n25603 = n10172 & n25602;
  assign n25604 = ~n8834 & n25603;
  assign n25605 = ~n9185 & n25604;
  assign n25606 = ~n9207 & n25605;
  assign n25607 = ~n9458 & n25606;
  assign n25608 = n9955 & n25607;
  assign n25609 = n9933 & n25608;
  assign n25610 = n10001 & n25609;
  assign n25611 = ~n25599 & ~n25610;
  assign n25612 = n25586 & n25611;
  assign n25613 = ~n8145 & n23844;
  assign n25614 = ~n9185 & n25613;
  assign n25615 = ~n9207 & n25614;
  assign n25616 = n9305 & n25615;
  assign n25617 = n9299 & n25616;
  assign n25618 = ~n7999 & n23894;
  assign n25619 = ~n9154 & n25618;
  assign n25620 = n9159 & n25619;
  assign n25621 = pi187 & ~n501;
  assign n25622 = n10133 & n25621;
  assign n25623 = n10138 & n25622;
  assign n25624 = n10131 & n25623;
  assign n25625 = ~n1172 & n25624;
  assign n25626 = ~n1114 & n25625;
  assign n25627 = ~n996 & n25626;
  assign n25628 = ~n500 & n25627;
  assign n25629 = n2316 & n25628;
  assign n25630 = n7608 & n25629;
  assign n25631 = n9915 & n25630;
  assign n25632 = n9856 & n25631;
  assign n25633 = n9733 & n25632;
  assign n25634 = ~n7236 & n25633;
  assign n25635 = ~n6137 & n25634;
  assign n25636 = n6193 & n25635;
  assign n25637 = n6134 & n25636;
  assign n25638 = ~n8867 & n25637;
  assign n25639 = ~n7235 & n25638;
  assign n25640 = n7296 & n25639;
  assign n25641 = n7231 & n25640;
  assign n25642 = ~n8866 & n25641;
  assign n25643 = n8898 & n25642;
  assign n25644 = n8863 & n25643;
  assign n25645 = ~n25620 & ~n25644;
  assign n25646 = ~n25617 & n25645;
  assign n25647 = ~n8053 & n23834;
  assign n25648 = ~n9185 & n25647;
  assign n25649 = ~n9206 & n25648;
  assign n25650 = n9214 & n25649;
  assign n25651 = ~n8218 & n23839;
  assign n25652 = ~n9185 & n25651;
  assign n25653 = n9324 & n25652;
  assign n25654 = n9379 & n25653;
  assign n25655 = n9373 & n25654;
  assign n25656 = ~n25650 & ~n25655;
  assign n25657 = n25646 & n25656;
  assign n25658 = n9282 & n21289;
  assign n25659 = ~n4817 & n25658;
  assign n25660 = ~n4902 & n25659;
  assign n25661 = ~n6001 & n25660;
  assign n25662 = ~n7014 & n25661;
  assign n25663 = ~n9261 & n25662;
  assign n25664 = ~n9185 & n25663;
  assign n25665 = ~n8114 & n25664;
  assign n25666 = ~n9260 & n25665;
  assign n25667 = n9259 & n25666;
  assign n25668 = n9253 & n25667;
  assign n25669 = n9246 & n25668;
  assign n25670 = n3846 & n22447;
  assign n25671 = n3854 & n25670;
  assign n25672 = n9138 & n25671;
  assign n25673 = ~n3066 & n25672;
  assign n25674 = ~n3983 & n25673;
  assign n25675 = ~n4003 & n25674;
  assign n25676 = ~n4024 & n25675;
  assign n25677 = ~n4999 & n25676;
  assign n25678 = ~n5827 & n25677;
  assign n25679 = ~n6893 & n25678;
  assign n25680 = ~n9114 & n25679;
  assign n25681 = ~n9113 & n25680;
  assign n25682 = ~n7890 & n25681;
  assign n25683 = ~n9112 & n25682;
  assign n25684 = n9111 & n25683;
  assign n25685 = n9104 & n25684;
  assign n25686 = n9097 & n25685;
  assign n25687 = ~n25669 & ~n25686;
  assign n25688 = n25657 & n25687;
  assign n25689 = n25612 & n25688;
  assign n25690 = n9355 & n21279;
  assign n25691 = ~n5808 & n25690;
  assign n25692 = ~n6056 & n25691;
  assign n25693 = ~n7073 & n25692;
  assign n25694 = ~n9330 & n25693;
  assign n25695 = ~n9185 & n25694;
  assign n25696 = ~n8179 & n25695;
  assign n25697 = ~n9329 & n25696;
  assign n25698 = n9328 & n25697;
  assign n25699 = n9323 & n25698;
  assign n25700 = n9316 & n25699;
  assign n25701 = ~n7204 & n23988;
  assign n25702 = ~n9185 & n25701;
  assign n25703 = ~n8291 & n25702;
  assign n25704 = ~n9444 & n25703;
  assign n25705 = n9450 & n25704;
  assign n25706 = n9443 & n25705;
  assign n25707 = n9442 & n25706;
  assign n25708 = ~n1208 & n23851;
  assign n25709 = n4920 & n25708;
  assign n25710 = ~n1270 & n25709;
  assign n25711 = n4932 & n25710;
  assign n25712 = ~n1372 & n25711;
  assign n25713 = ~n2243 & n25712;
  assign n25714 = ~n3104 & n25713;
  assign n25715 = ~n3971 & n25714;
  assign n25716 = ~n4003 & n25715;
  assign n25717 = ~n4872 & n25716;
  assign n25718 = ~n5801 & n25717;
  assign n25719 = ~n6739 & n25718;
  assign n25720 = ~n7807 & n25719;
  assign n25721 = ~n9070 & n25720;
  assign n25722 = ~n9069 & n25721;
  assign n25723 = ~n9068 & n25722;
  assign n25724 = ~n9067 & n25723;
  assign n25725 = n9066 & n25724;
  assign n25726 = n9060 & n25725;
  assign n25727 = n9053 & n25726;
  assign n25728 = ~n25707 & ~n25727;
  assign n25729 = ~n25700 & n25728;
  assign n25730 = n3740 & n19579;
  assign n25731 = n3951 & n25730;
  assign n25732 = n9220 & n25731;
  assign n25733 = ~n3940 & n25732;
  assign n25734 = ~n4001 & n25733;
  assign n25735 = ~n5043 & n25734;
  assign n25736 = ~n5943 & n25735;
  assign n25737 = ~n6951 & n25736;
  assign n25738 = ~n9186 & n25737;
  assign n25739 = ~n9185 & n25738;
  assign n25740 = ~n8037 & n25739;
  assign n25741 = ~n9184 & n25740;
  assign n25742 = n9183 & n25741;
  assign n25743 = n9176 & n25742;
  assign n25744 = n9169 & n25743;
  assign n25745 = pi163 & ~po161;
  assign n25746 = ~n9185 & n25745;
  assign n25747 = ~n8397 & n25746;
  assign n25748 = ~n9458 & n25747;
  assign n25749 = n9443 & n25748;
  assign n25750 = n10088 & n25749;
  assign n25751 = n10081 & n25750;
  assign n25752 = ~n25744 & ~n25751;
  assign n25753 = ~n1897 & n18618;
  assign n25754 = n1743 & n25753;
  assign n25755 = ~n2242 & n25754;
  assign n25756 = ~n3095 & n25755;
  assign n25757 = ~n3997 & n25756;
  assign n25758 = ~n4003 & n25757;
  assign n25759 = ~n4837 & n25758;
  assign n25760 = ~n5822 & n25759;
  assign n25761 = ~n6820 & n25760;
  assign n25762 = ~n7785 & n25761;
  assign n25763 = ~n9029 & n25762;
  assign n25764 = ~n9028 & n25763;
  assign n25765 = ~n9027 & n25764;
  assign n25766 = ~n9010 & n25765;
  assign n25767 = n9009 & n25766;
  assign n25768 = n9002 & n25767;
  assign n25769 = n8995 & n25768;
  assign n25770 = pi179 & ~n9511;
  assign n25771 = ~n8900 & n25770;
  assign n25772 = ~n9185 & n25771;
  assign n25773 = ~n9458 & n25772;
  assign n25774 = n9517 & n25773;
  assign n25775 = n9443 & n25774;
  assign n25776 = n9532 & n25775;
  assign n25777 = ~n25769 & ~n25776;
  assign n25778 = n25752 & n25777;
  assign n25779 = n25729 & n25778;
  assign po100 = ~n25689 | ~n25779;
  assign n25781 = pi196 & ~n501;
  assign n25782 = n5714 & n25781;
  assign n25783 = n5719 & n25782;
  assign n25784 = n8912 & n25783;
  assign n25785 = ~n1172 & n25784;
  assign n25786 = ~n996 & n25785;
  assign n25787 = ~n2306 & n25786;
  assign n25788 = ~n500 & n25787;
  assign n25789 = n2316 & n25788;
  assign n25790 = n7608 & n25789;
  assign n25791 = n10030 & n25790;
  assign n25792 = n10029 & n25791;
  assign n25793 = ~n7236 & n25792;
  assign n25794 = ~n6137 & n25793;
  assign n25795 = n6193 & n25794;
  assign n25796 = n6134 & n25795;
  assign n25797 = ~n8867 & n25796;
  assign n25798 = ~n7235 & n25797;
  assign n25799 = n7296 & n25798;
  assign n25800 = n7231 & n25799;
  assign n25801 = ~n10027 & n25800;
  assign n25802 = ~n8866 & n25801;
  assign n25803 = n8898 & n25802;
  assign n25804 = n8863 & n25803;
  assign n25805 = ~n10026 & n25804;
  assign n25806 = n10072 & n25805;
  assign n25807 = n10021 & n25806;
  assign n25808 = n8358 & n24206;
  assign n25809 = n9496 & n25808;
  assign n25810 = n9499 & n25809;
  assign n25811 = ~n7869 & n25810;
  assign n25812 = ~n9472 & n25811;
  assign n25813 = ~n9185 & n25812;
  assign n25814 = ~n8346 & n25813;
  assign n25815 = ~n9471 & n25814;
  assign n25816 = n9470 & n25815;
  assign n25817 = n9467 & n25816;
  assign n25818 = n9460 & n25817;
  assign n25819 = ~n25807 & ~n25818;
  assign n25820 = pi140 & ~n6461;
  assign n25821 = n6343 & n25820;
  assign n25822 = n8233 & n25821;
  assign n25823 = n9425 & n25822;
  assign n25824 = ~n6784 & n25823;
  assign n25825 = ~n7158 & n25824;
  assign n25826 = ~n9402 & n25825;
  assign n25827 = ~n9185 & n25826;
  assign n25828 = ~n8250 & n25827;
  assign n25829 = ~n9401 & n25828;
  assign n25830 = n9400 & n25829;
  assign n25831 = n9397 & n25830;
  assign n25832 = n9390 & n25831;
  assign n25833 = pi172 & ~n8762;
  assign n25834 = n8822 & n25833;
  assign n25835 = n8664 & n25834;
  assign n25836 = n10172 & n25835;
  assign n25837 = ~n8834 & n25836;
  assign n25838 = ~n9185 & n25837;
  assign n25839 = ~n9207 & n25838;
  assign n25840 = ~n9458 & n25839;
  assign n25841 = n9955 & n25840;
  assign n25842 = n9933 & n25841;
  assign n25843 = n10001 & n25842;
  assign n25844 = ~n25832 & ~n25843;
  assign n25845 = n25819 & n25844;
  assign n25846 = ~n8145 & n24049;
  assign n25847 = ~n9185 & n25846;
  assign n25848 = ~n9207 & n25847;
  assign n25849 = n9305 & n25848;
  assign n25850 = n9299 & n25849;
  assign n25851 = ~n7999 & n24078;
  assign n25852 = ~n9154 & n25851;
  assign n25853 = n9159 & n25852;
  assign n25854 = pi188 & ~n501;
  assign n25855 = n10133 & n25854;
  assign n25856 = n10138 & n25855;
  assign n25857 = n10131 & n25856;
  assign n25858 = ~n1172 & n25857;
  assign n25859 = ~n1114 & n25858;
  assign n25860 = ~n996 & n25859;
  assign n25861 = ~n500 & n25860;
  assign n25862 = n2316 & n25861;
  assign n25863 = n7608 & n25862;
  assign n25864 = n9915 & n25863;
  assign n25865 = n9856 & n25864;
  assign n25866 = n9733 & n25865;
  assign n25867 = ~n7236 & n25866;
  assign n25868 = ~n6137 & n25867;
  assign n25869 = n6193 & n25868;
  assign n25870 = n6134 & n25869;
  assign n25871 = ~n8867 & n25870;
  assign n25872 = ~n7235 & n25871;
  assign n25873 = n7296 & n25872;
  assign n25874 = n7231 & n25873;
  assign n25875 = ~n8866 & n25874;
  assign n25876 = n8898 & n25875;
  assign n25877 = n8863 & n25876;
  assign n25878 = ~n25853 & ~n25877;
  assign n25879 = ~n25850 & n25878;
  assign n25880 = ~n8053 & n24054;
  assign n25881 = ~n9185 & n25880;
  assign n25882 = ~n9206 & n25881;
  assign n25883 = n9214 & n25882;
  assign n25884 = ~n8218 & n24073;
  assign n25885 = ~n9185 & n25884;
  assign n25886 = n9324 & n25885;
  assign n25887 = n9379 & n25886;
  assign n25888 = n9373 & n25887;
  assign n25889 = ~n25883 & ~n25888;
  assign n25890 = n25879 & n25889;
  assign n25891 = n9282 & n21415;
  assign n25892 = ~n4817 & n25891;
  assign n25893 = ~n4902 & n25892;
  assign n25894 = ~n6001 & n25893;
  assign n25895 = ~n7014 & n25894;
  assign n25896 = ~n9261 & n25895;
  assign n25897 = ~n9185 & n25896;
  assign n25898 = ~n8114 & n25897;
  assign n25899 = ~n9260 & n25898;
  assign n25900 = n9259 & n25899;
  assign n25901 = n9253 & n25900;
  assign n25902 = n9246 & n25901;
  assign n25903 = n3846 & n22614;
  assign n25904 = n3854 & n25903;
  assign n25905 = n9138 & n25904;
  assign n25906 = ~n3066 & n25905;
  assign n25907 = ~n3983 & n25906;
  assign n25908 = ~n4003 & n25907;
  assign n25909 = ~n4024 & n25908;
  assign n25910 = ~n4999 & n25909;
  assign n25911 = ~n5827 & n25910;
  assign n25912 = ~n6893 & n25911;
  assign n25913 = ~n9114 & n25912;
  assign n25914 = ~n9113 & n25913;
  assign n25915 = ~n7890 & n25914;
  assign n25916 = ~n9112 & n25915;
  assign n25917 = n9111 & n25916;
  assign n25918 = n9104 & n25917;
  assign n25919 = n9097 & n25918;
  assign n25920 = ~n25902 & ~n25919;
  assign n25921 = n25890 & n25920;
  assign n25922 = n25845 & n25921;
  assign n25923 = n9355 & n21405;
  assign n25924 = ~n5808 & n25923;
  assign n25925 = ~n6056 & n25924;
  assign n25926 = ~n7073 & n25925;
  assign n25927 = ~n9330 & n25926;
  assign n25928 = ~n9185 & n25927;
  assign n25929 = ~n8179 & n25928;
  assign n25930 = ~n9329 & n25929;
  assign n25931 = n9328 & n25930;
  assign n25932 = n9323 & n25931;
  assign n25933 = n9316 & n25932;
  assign n25934 = ~n7204 & n24168;
  assign n25935 = ~n9185 & n25934;
  assign n25936 = ~n8291 & n25935;
  assign n25937 = ~n9444 & n25936;
  assign n25938 = n9450 & n25937;
  assign n25939 = n9443 & n25938;
  assign n25940 = n9442 & n25939;
  assign n25941 = ~n1208 & n24105;
  assign n25942 = n4920 & n25941;
  assign n25943 = ~n1270 & n25942;
  assign n25944 = n4932 & n25943;
  assign n25945 = ~n1372 & n25944;
  assign n25946 = ~n2243 & n25945;
  assign n25947 = ~n3104 & n25946;
  assign n25948 = ~n3971 & n25947;
  assign n25949 = ~n4003 & n25948;
  assign n25950 = ~n4872 & n25949;
  assign n25951 = ~n5801 & n25950;
  assign n25952 = ~n6739 & n25951;
  assign n25953 = ~n7807 & n25952;
  assign n25954 = ~n9070 & n25953;
  assign n25955 = ~n9069 & n25954;
  assign n25956 = ~n9068 & n25955;
  assign n25957 = ~n9067 & n25956;
  assign n25958 = n9066 & n25957;
  assign n25959 = n9060 & n25958;
  assign n25960 = n9053 & n25959;
  assign n25961 = ~n25940 & ~n25960;
  assign n25962 = ~n25933 & n25961;
  assign n25963 = n3740 & n19650;
  assign n25964 = n3951 & n25963;
  assign n25965 = n9220 & n25964;
  assign n25966 = ~n3940 & n25965;
  assign n25967 = ~n4001 & n25966;
  assign n25968 = ~n5043 & n25967;
  assign n25969 = ~n5943 & n25968;
  assign n25970 = ~n6951 & n25969;
  assign n25971 = ~n9186 & n25970;
  assign n25972 = ~n9185 & n25971;
  assign n25973 = ~n8037 & n25972;
  assign n25974 = ~n9184 & n25973;
  assign n25975 = n9183 & n25974;
  assign n25976 = n9176 & n25975;
  assign n25977 = n9169 & n25976;
  assign n25978 = pi164 & ~po161;
  assign n25979 = ~n9185 & n25978;
  assign n25980 = ~n8397 & n25979;
  assign n25981 = ~n9458 & n25980;
  assign n25982 = n9443 & n25981;
  assign n25983 = n10088 & n25982;
  assign n25984 = n10081 & n25983;
  assign n25985 = ~n25977 & ~n25984;
  assign n25986 = ~n1897 & n18656;
  assign n25987 = n1743 & n25986;
  assign n25988 = ~n2242 & n25987;
  assign n25989 = ~n3095 & n25988;
  assign n25990 = ~n3997 & n25989;
  assign n25991 = ~n4003 & n25990;
  assign n25992 = ~n4837 & n25991;
  assign n25993 = ~n5822 & n25992;
  assign n25994 = ~n6820 & n25993;
  assign n25995 = ~n7785 & n25994;
  assign n25996 = ~n9029 & n25995;
  assign n25997 = ~n9028 & n25996;
  assign n25998 = ~n9027 & n25997;
  assign n25999 = ~n9010 & n25998;
  assign n26000 = n9009 & n25999;
  assign n26001 = n9002 & n26000;
  assign n26002 = n8995 & n26001;
  assign n26003 = pi180 & ~n9511;
  assign n26004 = ~n8900 & n26003;
  assign n26005 = ~n9185 & n26004;
  assign n26006 = ~n9458 & n26005;
  assign n26007 = n9517 & n26006;
  assign n26008 = n9443 & n26007;
  assign n26009 = n9532 & n26008;
  assign n26010 = ~n26002 & ~n26009;
  assign n26011 = n25985 & n26010;
  assign n26012 = n25962 & n26011;
  assign po101 = ~n25922 | ~n26012;
  assign n26014 = pi197 & ~n501;
  assign n26015 = n5714 & n26014;
  assign n26016 = n5719 & n26015;
  assign n26017 = n8912 & n26016;
  assign n26018 = ~n1172 & n26017;
  assign n26019 = ~n996 & n26018;
  assign n26020 = ~n2306 & n26019;
  assign n26021 = ~n500 & n26020;
  assign n26022 = n2316 & n26021;
  assign n26023 = n7608 & n26022;
  assign n26024 = n10030 & n26023;
  assign n26025 = n10029 & n26024;
  assign n26026 = ~n7236 & n26025;
  assign n26027 = ~n6137 & n26026;
  assign n26028 = n6193 & n26027;
  assign n26029 = n6134 & n26028;
  assign n26030 = ~n8867 & n26029;
  assign n26031 = ~n7235 & n26030;
  assign n26032 = n7296 & n26031;
  assign n26033 = n7231 & n26032;
  assign n26034 = ~n10027 & n26033;
  assign n26035 = ~n8866 & n26034;
  assign n26036 = n8898 & n26035;
  assign n26037 = n8863 & n26036;
  assign n26038 = ~n10026 & n26037;
  assign n26039 = n10072 & n26038;
  assign n26040 = n10021 & n26039;
  assign n26041 = n8358 & n24399;
  assign n26042 = n9496 & n26041;
  assign n26043 = n9499 & n26042;
  assign n26044 = ~n7869 & n26043;
  assign n26045 = ~n9472 & n26044;
  assign n26046 = ~n9185 & n26045;
  assign n26047 = ~n8346 & n26046;
  assign n26048 = ~n9471 & n26047;
  assign n26049 = n9470 & n26048;
  assign n26050 = n9467 & n26049;
  assign n26051 = n9460 & n26050;
  assign n26052 = ~n26040 & ~n26051;
  assign n26053 = pi141 & ~n6461;
  assign n26054 = n6343 & n26053;
  assign n26055 = n8233 & n26054;
  assign n26056 = n9425 & n26055;
  assign n26057 = ~n6784 & n26056;
  assign n26058 = ~n7158 & n26057;
  assign n26059 = ~n9402 & n26058;
  assign n26060 = ~n9185 & n26059;
  assign n26061 = ~n8250 & n26060;
  assign n26062 = ~n9401 & n26061;
  assign n26063 = n9400 & n26062;
  assign n26064 = n9397 & n26063;
  assign n26065 = n9390 & n26064;
  assign n26066 = pi173 & ~n8762;
  assign n26067 = n8822 & n26066;
  assign n26068 = n8664 & n26067;
  assign n26069 = n10172 & n26068;
  assign n26070 = ~n8834 & n26069;
  assign n26071 = ~n9185 & n26070;
  assign n26072 = ~n9207 & n26071;
  assign n26073 = ~n9458 & n26072;
  assign n26074 = n9955 & n26073;
  assign n26075 = n9933 & n26074;
  assign n26076 = n10001 & n26075;
  assign n26077 = ~n26065 & ~n26076;
  assign n26078 = n26052 & n26077;
  assign n26079 = ~n8145 & n24242;
  assign n26080 = ~n9185 & n26079;
  assign n26081 = ~n9207 & n26080;
  assign n26082 = n9305 & n26081;
  assign n26083 = n9299 & n26082;
  assign n26084 = ~n7999 & n24271;
  assign n26085 = ~n9154 & n26084;
  assign n26086 = n9159 & n26085;
  assign n26087 = pi189 & ~n501;
  assign n26088 = n10133 & n26087;
  assign n26089 = n10138 & n26088;
  assign n26090 = n10131 & n26089;
  assign n26091 = ~n1172 & n26090;
  assign n26092 = ~n1114 & n26091;
  assign n26093 = ~n996 & n26092;
  assign n26094 = ~n500 & n26093;
  assign n26095 = n2316 & n26094;
  assign n26096 = n7608 & n26095;
  assign n26097 = n9915 & n26096;
  assign n26098 = n9856 & n26097;
  assign n26099 = n9733 & n26098;
  assign n26100 = ~n7236 & n26099;
  assign n26101 = ~n6137 & n26100;
  assign n26102 = n6193 & n26101;
  assign n26103 = n6134 & n26102;
  assign n26104 = ~n8867 & n26103;
  assign n26105 = ~n7235 & n26104;
  assign n26106 = n7296 & n26105;
  assign n26107 = n7231 & n26106;
  assign n26108 = ~n8866 & n26107;
  assign n26109 = n8898 & n26108;
  assign n26110 = n8863 & n26109;
  assign n26111 = ~n26086 & ~n26110;
  assign n26112 = ~n26083 & n26111;
  assign n26113 = ~n8053 & n24247;
  assign n26114 = ~n9185 & n26113;
  assign n26115 = ~n9206 & n26114;
  assign n26116 = n9214 & n26115;
  assign n26117 = ~n8218 & n24266;
  assign n26118 = ~n9185 & n26117;
  assign n26119 = n9324 & n26118;
  assign n26120 = n9379 & n26119;
  assign n26121 = n9373 & n26120;
  assign n26122 = ~n26116 & ~n26121;
  assign n26123 = n26112 & n26122;
  assign n26124 = n9282 & n21541;
  assign n26125 = ~n4817 & n26124;
  assign n26126 = ~n4902 & n26125;
  assign n26127 = ~n6001 & n26126;
  assign n26128 = ~n7014 & n26127;
  assign n26129 = ~n9261 & n26128;
  assign n26130 = ~n9185 & n26129;
  assign n26131 = ~n8114 & n26130;
  assign n26132 = ~n9260 & n26131;
  assign n26133 = n9259 & n26132;
  assign n26134 = n9253 & n26133;
  assign n26135 = n9246 & n26134;
  assign n26136 = n3846 & n22781;
  assign n26137 = n3854 & n26136;
  assign n26138 = n9138 & n26137;
  assign n26139 = ~n3066 & n26138;
  assign n26140 = ~n3983 & n26139;
  assign n26141 = ~n4003 & n26140;
  assign n26142 = ~n4024 & n26141;
  assign n26143 = ~n4999 & n26142;
  assign n26144 = ~n5827 & n26143;
  assign n26145 = ~n6893 & n26144;
  assign n26146 = ~n9114 & n26145;
  assign n26147 = ~n9113 & n26146;
  assign n26148 = ~n7890 & n26147;
  assign n26149 = ~n9112 & n26148;
  assign n26150 = n9111 & n26149;
  assign n26151 = n9104 & n26150;
  assign n26152 = n9097 & n26151;
  assign n26153 = ~n26135 & ~n26152;
  assign n26154 = n26123 & n26153;
  assign n26155 = n26078 & n26154;
  assign n26156 = n9355 & n21531;
  assign n26157 = ~n5808 & n26156;
  assign n26158 = ~n6056 & n26157;
  assign n26159 = ~n7073 & n26158;
  assign n26160 = ~n9330 & n26159;
  assign n26161 = ~n9185 & n26160;
  assign n26162 = ~n8179 & n26161;
  assign n26163 = ~n9329 & n26162;
  assign n26164 = n9328 & n26163;
  assign n26165 = n9323 & n26164;
  assign n26166 = n9316 & n26165;
  assign n26167 = ~n7204 & n24361;
  assign n26168 = ~n9185 & n26167;
  assign n26169 = ~n8291 & n26168;
  assign n26170 = ~n9444 & n26169;
  assign n26171 = n9450 & n26170;
  assign n26172 = n9443 & n26171;
  assign n26173 = n9442 & n26172;
  assign n26174 = ~n1208 & n24298;
  assign n26175 = n4920 & n26174;
  assign n26176 = ~n1270 & n26175;
  assign n26177 = n4932 & n26176;
  assign n26178 = ~n1372 & n26177;
  assign n26179 = ~n2243 & n26178;
  assign n26180 = ~n3104 & n26179;
  assign n26181 = ~n3971 & n26180;
  assign n26182 = ~n4003 & n26181;
  assign n26183 = ~n4872 & n26182;
  assign n26184 = ~n5801 & n26183;
  assign n26185 = ~n6739 & n26184;
  assign n26186 = ~n7807 & n26185;
  assign n26187 = ~n9070 & n26186;
  assign n26188 = ~n9069 & n26187;
  assign n26189 = ~n9068 & n26188;
  assign n26190 = ~n9067 & n26189;
  assign n26191 = n9066 & n26190;
  assign n26192 = n9060 & n26191;
  assign n26193 = n9053 & n26192;
  assign n26194 = ~n26173 & ~n26193;
  assign n26195 = ~n26166 & n26194;
  assign n26196 = n3740 & n19721;
  assign n26197 = n3951 & n26196;
  assign n26198 = n9220 & n26197;
  assign n26199 = ~n3940 & n26198;
  assign n26200 = ~n4001 & n26199;
  assign n26201 = ~n5043 & n26200;
  assign n26202 = ~n5943 & n26201;
  assign n26203 = ~n6951 & n26202;
  assign n26204 = ~n9186 & n26203;
  assign n26205 = ~n9185 & n26204;
  assign n26206 = ~n8037 & n26205;
  assign n26207 = ~n9184 & n26206;
  assign n26208 = n9183 & n26207;
  assign n26209 = n9176 & n26208;
  assign n26210 = n9169 & n26209;
  assign n26211 = pi165 & ~po161;
  assign n26212 = ~n9185 & n26211;
  assign n26213 = ~n8397 & n26212;
  assign n26214 = ~n9458 & n26213;
  assign n26215 = n9443 & n26214;
  assign n26216 = n10088 & n26215;
  assign n26217 = n10081 & n26216;
  assign n26218 = ~n26210 & ~n26217;
  assign n26219 = ~n1897 & n18694;
  assign n26220 = n1743 & n26219;
  assign n26221 = ~n2242 & n26220;
  assign n26222 = ~n3095 & n26221;
  assign n26223 = ~n3997 & n26222;
  assign n26224 = ~n4003 & n26223;
  assign n26225 = ~n4837 & n26224;
  assign n26226 = ~n5822 & n26225;
  assign n26227 = ~n6820 & n26226;
  assign n26228 = ~n7785 & n26227;
  assign n26229 = ~n9029 & n26228;
  assign n26230 = ~n9028 & n26229;
  assign n26231 = ~n9027 & n26230;
  assign n26232 = ~n9010 & n26231;
  assign n26233 = n9009 & n26232;
  assign n26234 = n9002 & n26233;
  assign n26235 = n8995 & n26234;
  assign n26236 = pi181 & ~n9511;
  assign n26237 = ~n8900 & n26236;
  assign n26238 = ~n9185 & n26237;
  assign n26239 = ~n9458 & n26238;
  assign n26240 = n9517 & n26239;
  assign n26241 = n9443 & n26240;
  assign n26242 = n9532 & n26241;
  assign n26243 = ~n26235 & ~n26242;
  assign n26244 = n26218 & n26243;
  assign n26245 = n26195 & n26244;
  assign po102 = ~n26155 | ~n26245;
  assign n26247 = pi198 & ~n501;
  assign n26248 = n5714 & n26247;
  assign n26249 = n5719 & n26248;
  assign n26250 = n8912 & n26249;
  assign n26251 = ~n1172 & n26250;
  assign n26252 = ~n996 & n26251;
  assign n26253 = ~n2306 & n26252;
  assign n26254 = ~n500 & n26253;
  assign n26255 = n2316 & n26254;
  assign n26256 = n7608 & n26255;
  assign n26257 = n10030 & n26256;
  assign n26258 = n10029 & n26257;
  assign n26259 = ~n7236 & n26258;
  assign n26260 = ~n6137 & n26259;
  assign n26261 = n6193 & n26260;
  assign n26262 = n6134 & n26261;
  assign n26263 = ~n8867 & n26262;
  assign n26264 = ~n7235 & n26263;
  assign n26265 = n7296 & n26264;
  assign n26266 = n7231 & n26265;
  assign n26267 = ~n10027 & n26266;
  assign n26268 = ~n8866 & n26267;
  assign n26269 = n8898 & n26268;
  assign n26270 = n8863 & n26269;
  assign n26271 = ~n10026 & n26270;
  assign n26272 = n10072 & n26271;
  assign n26273 = n10021 & n26272;
  assign n26274 = n8358 & n24592;
  assign n26275 = n9496 & n26274;
  assign n26276 = n9499 & n26275;
  assign n26277 = ~n7869 & n26276;
  assign n26278 = ~n9472 & n26277;
  assign n26279 = ~n9185 & n26278;
  assign n26280 = ~n8346 & n26279;
  assign n26281 = ~n9471 & n26280;
  assign n26282 = n9470 & n26281;
  assign n26283 = n9467 & n26282;
  assign n26284 = n9460 & n26283;
  assign n26285 = ~n26273 & ~n26284;
  assign n26286 = pi142 & ~n6461;
  assign n26287 = n6343 & n26286;
  assign n26288 = n8233 & n26287;
  assign n26289 = n9425 & n26288;
  assign n26290 = ~n6784 & n26289;
  assign n26291 = ~n7158 & n26290;
  assign n26292 = ~n9402 & n26291;
  assign n26293 = ~n9185 & n26292;
  assign n26294 = ~n8250 & n26293;
  assign n26295 = ~n9401 & n26294;
  assign n26296 = n9400 & n26295;
  assign n26297 = n9397 & n26296;
  assign n26298 = n9390 & n26297;
  assign n26299 = pi174 & ~n8762;
  assign n26300 = n8822 & n26299;
  assign n26301 = n8664 & n26300;
  assign n26302 = n10172 & n26301;
  assign n26303 = ~n8834 & n26302;
  assign n26304 = ~n9185 & n26303;
  assign n26305 = ~n9207 & n26304;
  assign n26306 = ~n9458 & n26305;
  assign n26307 = n9955 & n26306;
  assign n26308 = n9933 & n26307;
  assign n26309 = n10001 & n26308;
  assign n26310 = ~n26298 & ~n26309;
  assign n26311 = n26285 & n26310;
  assign n26312 = ~n8145 & n24435;
  assign n26313 = ~n9185 & n26312;
  assign n26314 = ~n9207 & n26313;
  assign n26315 = n9305 & n26314;
  assign n26316 = n9299 & n26315;
  assign n26317 = ~n7999 & n24464;
  assign n26318 = ~n9154 & n26317;
  assign n26319 = n9159 & n26318;
  assign n26320 = pi190 & ~n501;
  assign n26321 = n10133 & n26320;
  assign n26322 = n10138 & n26321;
  assign n26323 = n10131 & n26322;
  assign n26324 = ~n1172 & n26323;
  assign n26325 = ~n1114 & n26324;
  assign n26326 = ~n996 & n26325;
  assign n26327 = ~n500 & n26326;
  assign n26328 = n2316 & n26327;
  assign n26329 = n7608 & n26328;
  assign n26330 = n9915 & n26329;
  assign n26331 = n9856 & n26330;
  assign n26332 = n9733 & n26331;
  assign n26333 = ~n7236 & n26332;
  assign n26334 = ~n6137 & n26333;
  assign n26335 = n6193 & n26334;
  assign n26336 = n6134 & n26335;
  assign n26337 = ~n8867 & n26336;
  assign n26338 = ~n7235 & n26337;
  assign n26339 = n7296 & n26338;
  assign n26340 = n7231 & n26339;
  assign n26341 = ~n8866 & n26340;
  assign n26342 = n8898 & n26341;
  assign n26343 = n8863 & n26342;
  assign n26344 = ~n26319 & ~n26343;
  assign n26345 = ~n26316 & n26344;
  assign n26346 = ~n8053 & n24440;
  assign n26347 = ~n9185 & n26346;
  assign n26348 = ~n9206 & n26347;
  assign n26349 = n9214 & n26348;
  assign n26350 = ~n8218 & n24459;
  assign n26351 = ~n9185 & n26350;
  assign n26352 = n9324 & n26351;
  assign n26353 = n9379 & n26352;
  assign n26354 = n9373 & n26353;
  assign n26355 = ~n26349 & ~n26354;
  assign n26356 = n26345 & n26355;
  assign n26357 = n9282 & n21667;
  assign n26358 = ~n4817 & n26357;
  assign n26359 = ~n4902 & n26358;
  assign n26360 = ~n6001 & n26359;
  assign n26361 = ~n7014 & n26360;
  assign n26362 = ~n9261 & n26361;
  assign n26363 = ~n9185 & n26362;
  assign n26364 = ~n8114 & n26363;
  assign n26365 = ~n9260 & n26364;
  assign n26366 = n9259 & n26365;
  assign n26367 = n9253 & n26366;
  assign n26368 = n9246 & n26367;
  assign n26369 = n3846 & n22948;
  assign n26370 = n3854 & n26369;
  assign n26371 = n9138 & n26370;
  assign n26372 = ~n3066 & n26371;
  assign n26373 = ~n3983 & n26372;
  assign n26374 = ~n4003 & n26373;
  assign n26375 = ~n4024 & n26374;
  assign n26376 = ~n4999 & n26375;
  assign n26377 = ~n5827 & n26376;
  assign n26378 = ~n6893 & n26377;
  assign n26379 = ~n9114 & n26378;
  assign n26380 = ~n9113 & n26379;
  assign n26381 = ~n7890 & n26380;
  assign n26382 = ~n9112 & n26381;
  assign n26383 = n9111 & n26382;
  assign n26384 = n9104 & n26383;
  assign n26385 = n9097 & n26384;
  assign n26386 = ~n26368 & ~n26385;
  assign n26387 = n26356 & n26386;
  assign n26388 = n26311 & n26387;
  assign n26389 = n9355 & n21657;
  assign n26390 = ~n5808 & n26389;
  assign n26391 = ~n6056 & n26390;
  assign n26392 = ~n7073 & n26391;
  assign n26393 = ~n9330 & n26392;
  assign n26394 = ~n9185 & n26393;
  assign n26395 = ~n8179 & n26394;
  assign n26396 = ~n9329 & n26395;
  assign n26397 = n9328 & n26396;
  assign n26398 = n9323 & n26397;
  assign n26399 = n9316 & n26398;
  assign n26400 = ~n7204 & n24554;
  assign n26401 = ~n9185 & n26400;
  assign n26402 = ~n8291 & n26401;
  assign n26403 = ~n9444 & n26402;
  assign n26404 = n9450 & n26403;
  assign n26405 = n9443 & n26404;
  assign n26406 = n9442 & n26405;
  assign n26407 = ~n1208 & n24491;
  assign n26408 = n4920 & n26407;
  assign n26409 = ~n1270 & n26408;
  assign n26410 = n4932 & n26409;
  assign n26411 = ~n1372 & n26410;
  assign n26412 = ~n2243 & n26411;
  assign n26413 = ~n3104 & n26412;
  assign n26414 = ~n3971 & n26413;
  assign n26415 = ~n4003 & n26414;
  assign n26416 = ~n4872 & n26415;
  assign n26417 = ~n5801 & n26416;
  assign n26418 = ~n6739 & n26417;
  assign n26419 = ~n7807 & n26418;
  assign n26420 = ~n9070 & n26419;
  assign n26421 = ~n9069 & n26420;
  assign n26422 = ~n9068 & n26421;
  assign n26423 = ~n9067 & n26422;
  assign n26424 = n9066 & n26423;
  assign n26425 = n9060 & n26424;
  assign n26426 = n9053 & n26425;
  assign n26427 = ~n26406 & ~n26426;
  assign n26428 = ~n26399 & n26427;
  assign n26429 = n3740 & n19792;
  assign n26430 = n3951 & n26429;
  assign n26431 = n9220 & n26430;
  assign n26432 = ~n3940 & n26431;
  assign n26433 = ~n4001 & n26432;
  assign n26434 = ~n5043 & n26433;
  assign n26435 = ~n5943 & n26434;
  assign n26436 = ~n6951 & n26435;
  assign n26437 = ~n9186 & n26436;
  assign n26438 = ~n9185 & n26437;
  assign n26439 = ~n8037 & n26438;
  assign n26440 = ~n9184 & n26439;
  assign n26441 = n9183 & n26440;
  assign n26442 = n9176 & n26441;
  assign n26443 = n9169 & n26442;
  assign n26444 = pi166 & ~po161;
  assign n26445 = ~n9185 & n26444;
  assign n26446 = ~n8397 & n26445;
  assign n26447 = ~n9458 & n26446;
  assign n26448 = n9443 & n26447;
  assign n26449 = n10088 & n26448;
  assign n26450 = n10081 & n26449;
  assign n26451 = ~n26443 & ~n26450;
  assign n26452 = ~n1897 & n18732;
  assign n26453 = n1743 & n26452;
  assign n26454 = ~n2242 & n26453;
  assign n26455 = ~n3095 & n26454;
  assign n26456 = ~n3997 & n26455;
  assign n26457 = ~n4003 & n26456;
  assign n26458 = ~n4837 & n26457;
  assign n26459 = ~n5822 & n26458;
  assign n26460 = ~n6820 & n26459;
  assign n26461 = ~n7785 & n26460;
  assign n26462 = ~n9029 & n26461;
  assign n26463 = ~n9028 & n26462;
  assign n26464 = ~n9027 & n26463;
  assign n26465 = ~n9010 & n26464;
  assign n26466 = n9009 & n26465;
  assign n26467 = n9002 & n26466;
  assign n26468 = n8995 & n26467;
  assign n26469 = pi182 & ~n9511;
  assign n26470 = ~n8900 & n26469;
  assign n26471 = ~n9185 & n26470;
  assign n26472 = ~n9458 & n26471;
  assign n26473 = n9517 & n26472;
  assign n26474 = n9443 & n26473;
  assign n26475 = n9532 & n26474;
  assign n26476 = ~n26468 & ~n26475;
  assign n26477 = n26451 & n26476;
  assign n26478 = n26428 & n26477;
  assign po103 = ~n26388 | ~n26478;
  assign n26480 = n11274 & n24609;
  assign n26481 = n8545 & n26480;
  assign n26482 = ~n8834 & n26481;
  assign n26483 = ~n11273 & n26482;
  assign n26484 = ~n10416 & n26483;
  assign n26485 = ~n10002 & n26484;
  assign n26486 = ~n10780 & n26485;
  assign n26487 = n10640 & n26486;
  assign n26488 = n11272 & n26487;
  assign n26489 = n11296 & n26488;
  assign n26490 = pi191 & ~n11324;
  assign n26491 = ~n10416 & n26490;
  assign n26492 = ~n10074 & n26491;
  assign n26493 = ~n10780 & n26492;
  assign n26494 = n10640 & n26493;
  assign n26495 = n11323 & n26494;
  assign n26496 = n11342 & n26495;
  assign n26497 = ~n26489 & ~n26496;
  assign n26498 = n8362 & n8364;
  assign n26499 = n8360 & n24742;
  assign n26500 = n26498 & n26499;
  assign n26501 = ~n7869 & n26500;
  assign n26502 = ~n8346 & n26501;
  assign n26503 = ~n10714 & n26502;
  assign n26504 = ~n10416 & n26503;
  assign n26505 = ~n9485 & n26504;
  assign n26506 = ~n10713 & n26505;
  assign n26507 = n10640 & n26506;
  assign n26508 = n10712 & n26507;
  assign n26509 = n10740 & n26508;
  assign n26510 = ~n4341 & ~n4489;
  assign n26511 = n4609 & n26510;
  assign n26512 = pi103 & ~n4307;
  assign n26513 = ~n4308 & n26512;
  assign n26514 = ~n4306 & n26513;
  assign n26515 = ~n4707 & n26514;
  assign n26516 = n5085 & n26515;
  assign n26517 = n26511 & n26516;
  assign n26518 = ~n4817 & n26517;
  assign n26519 = ~n4902 & n26518;
  assign n26520 = ~n6001 & n26519;
  assign n26521 = ~n7014 & n26520;
  assign n26522 = ~n8114 & n26521;
  assign n26523 = ~n10496 & n26522;
  assign n26524 = ~n10416 & n26523;
  assign n26525 = ~n9276 & n26524;
  assign n26526 = ~n10495 & n26525;
  assign n26527 = n10494 & n26526;
  assign n26528 = n10490 & n26527;
  assign n26529 = n10522 & n26528;
  assign n26530 = ~n26509 & ~n26529;
  assign n26531 = n26497 & n26530;
  assign n26532 = ~n9215 & n24701;
  assign n26533 = ~n10416 & n26532;
  assign n26534 = ~n10451 & n26533;
  assign n26535 = n10459 & n26534;
  assign n26536 = ~n9160 & n24691;
  assign n26537 = ~n10394 & n26536;
  assign n26538 = n10399 & n26537;
  assign n26539 = pi199 & ~n501;
  assign n26540 = n11440 & n26539;
  assign n26541 = n11446 & n26540;
  assign n26542 = n11437 & n26541;
  assign n26543 = ~n1172 & n26542;
  assign n26544 = ~n996 & n26543;
  assign n26545 = ~n2306 & n26544;
  assign n26546 = ~n500 & n26545;
  assign n26547 = n11004 & n26546;
  assign n26548 = ~n2482 & ~n3254;
  assign n26549 = n11006 & n26548;
  assign n26550 = n21846 & n26549;
  assign n26551 = n26547 & n26550;
  assign n26552 = n10980 & n26551;
  assign n26553 = n10971 & n26552;
  assign n26554 = n11172 & n26553;
  assign n26555 = ~n7236 & n26554;
  assign n26556 = ~n6137 & n26555;
  assign n26557 = n6193 & n26556;
  assign n26558 = n6134 & n26557;
  assign n26559 = ~n8867 & n26558;
  assign n26560 = ~n7235 & n26559;
  assign n26561 = n7296 & n26560;
  assign n26562 = n7231 & n26561;
  assign n26563 = ~n10027 & n26562;
  assign n26564 = ~n8866 & n26563;
  assign n26565 = n8898 & n26564;
  assign n26566 = n8863 & n26565;
  assign n26567 = ~n10026 & n26566;
  assign n26568 = n10072 & n26567;
  assign n26569 = n10021 & n26568;
  assign n26570 = pi207 & ~n501;
  assign n26571 = n4792 & n12872;
  assign n26572 = n26570 & n26571;
  assign n26573 = n14210 & n15998;
  assign n26574 = n12604 & n26573;
  assign n26575 = n11411 & n26574;
  assign n26576 = n26572 & n26575;
  assign n26577 = n11404 & n26576;
  assign n26578 = ~n1172 & n26577;
  assign n26579 = ~n996 & n26578;
  assign n26580 = ~n2306 & n26579;
  assign n26581 = ~n500 & n26580;
  assign n26582 = n10855 & n26581;
  assign n26583 = n10857 & n12578;
  assign n26584 = n21846 & n26583;
  assign n26585 = n26582 & n26584;
  assign n26586 = n10831 & n26585;
  assign n26587 = n10823 & n26586;
  assign n26588 = ~n7236 & n26587;
  assign n26589 = ~n6137 & n26588;
  assign n26590 = n6193 & n26589;
  assign n26591 = n6134 & n26590;
  assign n26592 = ~n8867 & n26591;
  assign n26593 = ~n7235 & n26592;
  assign n26594 = n7296 & n26593;
  assign n26595 = n7231 & n26594;
  assign n26596 = ~n10027 & n26595;
  assign n26597 = ~n8866 & n26596;
  assign n26598 = n8898 & n26597;
  assign n26599 = n8863 & n26598;
  assign n26600 = ~n10788 & n26599;
  assign n26601 = ~n10026 & n26600;
  assign n26602 = n10072 & n26601;
  assign n26603 = n10021 & n26602;
  assign n26604 = ~n26569 & ~n26603;
  assign n26605 = ~n26538 & n26604;
  assign n26606 = ~n26535 & n26605;
  assign n26607 = ~n9381 & n24662;
  assign n26608 = ~n10416 & n26607;
  assign n26609 = n10564 & n26608;
  assign n26610 = n10627 & n26609;
  assign n26611 = n10621 & n26610;
  assign n26612 = ~n9307 & n24696;
  assign n26613 = ~n10416 & n26612;
  assign n26614 = ~n10452 & n26613;
  assign n26615 = n10552 & n26614;
  assign n26616 = n10546 & n26615;
  assign n26617 = ~n26611 & ~n26616;
  assign n26618 = n26606 & n26617;
  assign n26619 = pi119 & ~n5598;
  assign n26620 = n6068 & n26619;
  assign n26621 = n6066 & n26620;
  assign n26622 = n10602 & n26621;
  assign n26623 = ~n5808 & n26622;
  assign n26624 = ~n6056 & n26623;
  assign n26625 = ~n7073 & n26624;
  assign n26626 = ~n8179 & n26625;
  assign n26627 = ~n10568 & n26626;
  assign n26628 = ~n10416 & n26627;
  assign n26629 = ~n9344 & n26628;
  assign n26630 = ~n10567 & n26629;
  assign n26631 = n10566 & n26630;
  assign n26632 = n10563 & n26631;
  assign n26633 = n10593 & n26632;
  assign n26634 = n9794 & ~n9824;
  assign n26635 = pi183 & pi255;
  assign n26636 = ~n9850 & n26635;
  assign n26637 = ~n9687 & n26636;
  assign n26638 = ~n9913 & n26637;
  assign n26639 = n11365 & n26638;
  assign n26640 = n26634 & n26639;
  assign n26641 = ~n9929 & n26640;
  assign n26642 = ~n10416 & n26641;
  assign n26643 = ~n10622 & n26642;
  assign n26644 = n10564 & n26643;
  assign n26645 = n11226 & n26644;
  assign n26646 = n11218 & n26645;
  assign n26647 = n11265 & n26646;
  assign n26648 = ~n26633 & ~n26647;
  assign n26649 = n26618 & n26648;
  assign n26650 = n26531 & n26649;
  assign n26651 = pi175 & ~n8900;
  assign n26652 = ~n10416 & n26651;
  assign n26653 = ~n9533 & n26652;
  assign n26654 = ~n10764 & n26653;
  assign n26655 = n10770 & n26654;
  assign n26656 = n10640 & n26655;
  assign n26657 = n10786 & n26656;
  assign n26658 = ~n8291 & n24653;
  assign n26659 = ~n10416 & n26658;
  assign n26660 = ~n9453 & n26659;
  assign n26661 = ~n10696 & n26660;
  assign n26662 = n10702 & n26661;
  assign n26663 = n10640 & n26662;
  assign n26664 = n10695 & n26663;
  assign n26665 = ~n26657 & ~n26664;
  assign n26666 = ~n8397 & n24714;
  assign n26667 = ~n10416 & n26666;
  assign n26668 = ~n10094 & n26667;
  assign n26669 = ~n10713 & n26668;
  assign n26670 = n10640 & n26669;
  assign n26671 = n11312 & n26670;
  assign n26672 = n11305 & n26671;
  assign n26673 = n5008 & n21712;
  assign n26674 = ~n3066 & n26673;
  assign n26675 = ~n3983 & n26674;
  assign n26676 = ~n4003 & n26675;
  assign n26677 = ~n4024 & n26676;
  assign n26678 = ~n4999 & n26677;
  assign n26679 = ~n5827 & n26678;
  assign n26680 = ~n6893 & n26679;
  assign n26681 = ~n7890 & n26680;
  assign n26682 = ~n10206 & n26681;
  assign n26683 = ~n10205 & n26682;
  assign n26684 = ~n9131 & n26683;
  assign n26685 = ~n10204 & n26684;
  assign n26686 = n10203 & n26685;
  assign n26687 = n10198 & n26686;
  assign n26688 = n10277 & n26687;
  assign n26689 = ~n26672 & ~n26688;
  assign n26690 = n26665 & n26689;
  assign n26691 = n719 & n4930;
  assign n26692 = pi039 & ~n653;
  assign n26693 = ~n654 & n26692;
  assign n26694 = ~n652 & n26693;
  assign n26695 = ~n1208 & n26694;
  assign n26696 = n11681 & n26695;
  assign n26697 = n26691 & n26696;
  assign n26698 = ~n1372 & n26697;
  assign n26699 = ~n2243 & n26698;
  assign n26700 = ~n3104 & n26699;
  assign n26701 = ~n3971 & n26700;
  assign n26702 = ~n4003 & n26701;
  assign n26703 = ~n4872 & n26702;
  assign n26704 = ~n5801 & n26703;
  assign n26705 = ~n6739 & n26704;
  assign n26706 = ~n7807 & n26705;
  assign n26707 = ~n8989 & n26706;
  assign n26708 = ~n10293 & n26707;
  assign n26709 = ~n10292 & n26708;
  assign n26710 = ~n10273 & n26709;
  assign n26711 = ~n10291 & n26710;
  assign n26712 = n10290 & n26711;
  assign n26713 = n10285 & n26712;
  assign n26714 = n10326 & n26713;
  assign n26715 = n4100 & n4103;
  assign n26716 = ~n3710 & n20681;
  assign n26717 = n5062 & n26716;
  assign n26718 = n26715 & n26717;
  assign n26719 = ~n3940 & n26718;
  assign n26720 = ~n4001 & n26719;
  assign n26721 = ~n5043 & n26720;
  assign n26722 = ~n5943 & n26721;
  assign n26723 = ~n6951 & n26722;
  assign n26724 = ~n8037 & n26723;
  assign n26725 = ~n10417 & n26724;
  assign n26726 = ~n10416 & n26725;
  assign n26727 = ~n9200 & n26726;
  assign n26728 = ~n10415 & n26727;
  assign n26729 = n10414 & n26728;
  assign n26730 = n10409 & n26729;
  assign n26731 = n10444 & n26730;
  assign n26732 = ~n26714 & ~n26731;
  assign n26733 = n6523 & n7176;
  assign n26734 = pi135 & ~n6668;
  assign n26735 = ~n6669 & n26734;
  assign n26736 = ~n6667 & n26735;
  assign n26737 = ~n6313 & n26736;
  assign n26738 = n7169 & n7175;
  assign n26739 = n26737 & n26738;
  assign n26740 = n26733 & n26739;
  assign n26741 = ~n6784 & n26740;
  assign n26742 = ~n7158 & n26741;
  assign n26743 = ~n8250 & n26742;
  assign n26744 = ~n10642 & n26743;
  assign n26745 = ~n10416 & n26744;
  assign n26746 = ~n9414 & n26745;
  assign n26747 = ~n10641 & n26746;
  assign n26748 = n10640 & n26747;
  assign n26749 = n10638 & n26748;
  assign n26750 = n10666 & n26749;
  assign n26751 = pi055 & ~n2139;
  assign n26752 = ~n2140 & n26751;
  assign n26753 = ~n2138 & n26752;
  assign n26754 = ~n2176 & n26753;
  assign n26755 = n11518 & n26754;
  assign n26756 = n1619 & n26755;
  assign n26757 = ~n2242 & n26756;
  assign n26758 = ~n3095 & n26757;
  assign n26759 = ~n3997 & n26758;
  assign n26760 = ~n4003 & n26759;
  assign n26761 = ~n4837 & n26760;
  assign n26762 = ~n5822 & n26761;
  assign n26763 = ~n6820 & n26762;
  assign n26764 = ~n7785 & n26763;
  assign n26765 = ~n9027 & n26764;
  assign n26766 = ~n10342 & n26765;
  assign n26767 = ~n10341 & n26766;
  assign n26768 = ~n10245 & n26767;
  assign n26769 = ~n10340 & n26768;
  assign n26770 = n10339 & n26769;
  assign n26771 = n10334 & n26770;
  assign n26772 = n10372 & n26771;
  assign n26773 = ~n26750 & ~n26772;
  assign n26774 = n26732 & n26773;
  assign n26775 = n26690 & n26774;
  assign po104 = ~n26650 | ~n26775;
  assign n26777 = n8363 & n24850;
  assign n26778 = ~n7869 & n26777;
  assign n26779 = ~n8346 & n26778;
  assign n26780 = ~n10714 & n26779;
  assign n26781 = ~n10416 & n26780;
  assign n26782 = ~n9485 & n26781;
  assign n26783 = ~n10713 & n26782;
  assign n26784 = n10640 & n26783;
  assign n26785 = n10712 & n26784;
  assign n26786 = n10740 & n26785;
  assign n26787 = pi088 & ~n3710;
  assign n26788 = n4096 & n26787;
  assign n26789 = n4104 & n26788;
  assign n26790 = n8056 & n26789;
  assign n26791 = ~n3940 & n26790;
  assign n26792 = ~n4001 & n26791;
  assign n26793 = ~n5043 & n26792;
  assign n26794 = ~n5943 & n26793;
  assign n26795 = ~n6951 & n26794;
  assign n26796 = ~n8037 & n26795;
  assign n26797 = ~n10417 & n26796;
  assign n26798 = ~n10416 & n26797;
  assign n26799 = ~n9200 & n26798;
  assign n26800 = ~n10415 & n26799;
  assign n26801 = n10414 & n26800;
  assign n26802 = n10409 & n26801;
  assign n26803 = n10444 & n26802;
  assign n26804 = ~n26786 & ~n26803;
  assign n26805 = n11378 & n24971;
  assign n26806 = n9942 & n26805;
  assign n26807 = ~n8834 & n26806;
  assign n26808 = ~n11273 & n26807;
  assign n26809 = ~n10416 & n26808;
  assign n26810 = ~n10002 & n26809;
  assign n26811 = ~n10780 & n26810;
  assign n26812 = n10640 & n26811;
  assign n26813 = n11272 & n26812;
  assign n26814 = n11296 & n26813;
  assign n26815 = pi104 & ~n4707;
  assign n26816 = n5083 & n26815;
  assign n26817 = n8096 & n26816;
  assign n26818 = n9263 & n26817;
  assign n26819 = ~n4817 & n26818;
  assign n26820 = ~n4902 & n26819;
  assign n26821 = ~n6001 & n26820;
  assign n26822 = ~n7014 & n26821;
  assign n26823 = ~n8114 & n26822;
  assign n26824 = ~n10496 & n26823;
  assign n26825 = ~n10416 & n26824;
  assign n26826 = ~n9276 & n26825;
  assign n26827 = ~n10495 & n26826;
  assign n26828 = n10494 & n26827;
  assign n26829 = n10490 & n26828;
  assign n26830 = n10522 & n26829;
  assign n26831 = ~n26814 & ~n26830;
  assign n26832 = n26804 & n26831;
  assign n26833 = ~n9215 & n24913;
  assign n26834 = ~n10416 & n26833;
  assign n26835 = ~n10451 & n26834;
  assign n26836 = n10459 & n26835;
  assign n26837 = ~n9160 & n24941;
  assign n26838 = ~n10394 & n26837;
  assign n26839 = n10399 & n26838;
  assign n26840 = pi200 & ~n501;
  assign n26841 = n11440 & n26840;
  assign n26842 = n11446 & n26841;
  assign n26843 = n11437 & n26842;
  assign n26844 = ~n1172 & n26843;
  assign n26845 = ~n996 & n26844;
  assign n26846 = ~n2306 & n26845;
  assign n26847 = ~n500 & n26846;
  assign n26848 = n11004 & n26847;
  assign n26849 = n26550 & n26848;
  assign n26850 = n10980 & n26849;
  assign n26851 = n10971 & n26850;
  assign n26852 = n11172 & n26851;
  assign n26853 = ~n7236 & n26852;
  assign n26854 = ~n6137 & n26853;
  assign n26855 = n6193 & n26854;
  assign n26856 = n6134 & n26855;
  assign n26857 = ~n8867 & n26856;
  assign n26858 = ~n7235 & n26857;
  assign n26859 = n7296 & n26858;
  assign n26860 = n7231 & n26859;
  assign n26861 = ~n10027 & n26860;
  assign n26862 = ~n8866 & n26861;
  assign n26863 = n8898 & n26862;
  assign n26864 = n8863 & n26863;
  assign n26865 = ~n10026 & n26864;
  assign n26866 = n10072 & n26865;
  assign n26867 = n10021 & n26866;
  assign n26868 = pi208 & ~n501;
  assign n26869 = n26571 & n26868;
  assign n26870 = n26575 & n26869;
  assign n26871 = n11404 & n26870;
  assign n26872 = ~n1172 & n26871;
  assign n26873 = ~n996 & n26872;
  assign n26874 = ~n2306 & n26873;
  assign n26875 = ~n500 & n26874;
  assign n26876 = n10855 & n26875;
  assign n26877 = n26584 & n26876;
  assign n26878 = n10831 & n26877;
  assign n26879 = n10823 & n26878;
  assign n26880 = ~n7236 & n26879;
  assign n26881 = ~n6137 & n26880;
  assign n26882 = n6193 & n26881;
  assign n26883 = n6134 & n26882;
  assign n26884 = ~n8867 & n26883;
  assign n26885 = ~n7235 & n26884;
  assign n26886 = n7296 & n26885;
  assign n26887 = n7231 & n26886;
  assign n26888 = ~n10027 & n26887;
  assign n26889 = ~n8866 & n26888;
  assign n26890 = n8898 & n26889;
  assign n26891 = n8863 & n26890;
  assign n26892 = ~n10788 & n26891;
  assign n26893 = ~n10026 & n26892;
  assign n26894 = n10072 & n26893;
  assign n26895 = n10021 & n26894;
  assign n26896 = ~n26867 & ~n26895;
  assign n26897 = ~n26839 & n26896;
  assign n26898 = ~n26836 & n26897;
  assign n26899 = ~n9307 & n24946;
  assign n26900 = ~n10416 & n26899;
  assign n26901 = ~n10452 & n26900;
  assign n26902 = n10552 & n26901;
  assign n26903 = n10546 & n26902;
  assign n26904 = ~n9381 & n24951;
  assign n26905 = ~n10416 & n26904;
  assign n26906 = n10564 & n26905;
  assign n26907 = n10627 & n26906;
  assign n26908 = n10621 & n26907;
  assign n26909 = ~n26903 & ~n26908;
  assign n26910 = n26898 & n26909;
  assign n26911 = n10602 & n20901;
  assign n26912 = ~n5808 & n26911;
  assign n26913 = ~n6056 & n26912;
  assign n26914 = ~n7073 & n26913;
  assign n26915 = ~n8179 & n26914;
  assign n26916 = ~n10568 & n26915;
  assign n26917 = ~n10416 & n26916;
  assign n26918 = ~n9344 & n26917;
  assign n26919 = ~n10567 & n26918;
  assign n26920 = n10566 & n26919;
  assign n26921 = n10563 & n26920;
  assign n26922 = n10593 & n26921;
  assign n26923 = pi184 & ~n9687;
  assign n26924 = ~n9913 & n26923;
  assign n26925 = n11365 & n26924;
  assign n26926 = n9856 & n26925;
  assign n26927 = ~n9929 & n26926;
  assign n26928 = ~n10416 & n26927;
  assign n26929 = ~n10622 & n26928;
  assign n26930 = n10564 & n26929;
  assign n26931 = n11226 & n26930;
  assign n26932 = n11218 & n26931;
  assign n26933 = n11265 & n26932;
  assign n26934 = ~n26922 & ~n26933;
  assign n26935 = n26910 & n26934;
  assign n26936 = n26832 & n26935;
  assign n26937 = pi192 & ~n11324;
  assign n26938 = ~n10416 & n26937;
  assign n26939 = ~n10074 & n26938;
  assign n26940 = ~n10780 & n26939;
  assign n26941 = n10640 & n26940;
  assign n26942 = n11323 & n26941;
  assign n26943 = n11342 & n26942;
  assign n26944 = pi176 & ~n8900;
  assign n26945 = ~n10416 & n26944;
  assign n26946 = ~n9533 & n26945;
  assign n26947 = ~n10764 & n26946;
  assign n26948 = n10770 & n26947;
  assign n26949 = n10640 & n26948;
  assign n26950 = n10786 & n26949;
  assign n26951 = ~n26943 & ~n26950;
  assign n26952 = pi040 & ~n1208;
  assign n26953 = n4920 & n26952;
  assign n26954 = n4931 & n26953;
  assign n26955 = n4928 & n26954;
  assign n26956 = ~n1372 & n26955;
  assign n26957 = ~n2243 & n26956;
  assign n26958 = ~n3104 & n26957;
  assign n26959 = ~n3971 & n26958;
  assign n26960 = ~n4003 & n26959;
  assign n26961 = ~n4872 & n26960;
  assign n26962 = ~n5801 & n26961;
  assign n26963 = ~n6739 & n26962;
  assign n26964 = ~n7807 & n26963;
  assign n26965 = ~n8989 & n26964;
  assign n26966 = ~n10293 & n26965;
  assign n26967 = ~n10292 & n26966;
  assign n26968 = ~n10273 & n26967;
  assign n26969 = ~n10291 & n26968;
  assign n26970 = n10290 & n26969;
  assign n26971 = n10285 & n26970;
  assign n26972 = n10326 & n26971;
  assign n26973 = ~n8397 & n24999;
  assign n26974 = ~n10416 & n26973;
  assign n26975 = ~n10094 & n26974;
  assign n26976 = ~n10713 & n26975;
  assign n26977 = n10640 & n26976;
  assign n26978 = n11312 & n26977;
  assign n26979 = n11305 & n26978;
  assign n26980 = ~n26972 & ~n26979;
  assign n26981 = n26951 & n26980;
  assign n26982 = ~n8291 & n25060;
  assign n26983 = ~n10416 & n26982;
  assign n26984 = ~n9453 & n26983;
  assign n26985 = ~n10696 & n26984;
  assign n26986 = n10702 & n26985;
  assign n26987 = n10640 & n26986;
  assign n26988 = n10695 & n26987;
  assign n26989 = n10376 & n24860;
  assign n26990 = n9115 & n26989;
  assign n26991 = ~n3066 & n26990;
  assign n26992 = ~n3983 & n26991;
  assign n26993 = ~n4003 & n26992;
  assign n26994 = ~n4024 & n26993;
  assign n26995 = ~n4999 & n26994;
  assign n26996 = ~n5827 & n26995;
  assign n26997 = ~n6893 & n26996;
  assign n26998 = ~n7890 & n26997;
  assign n26999 = ~n10206 & n26998;
  assign n27000 = ~n10205 & n26999;
  assign n27001 = ~n9131 & n27000;
  assign n27002 = ~n10204 & n27001;
  assign n27003 = n10203 & n27002;
  assign n27004 = n10198 & n27003;
  assign n27005 = n10277 & n27004;
  assign n27006 = ~n26988 & ~n27005;
  assign n27007 = pi136 & ~n6313;
  assign n27008 = n7169 & n27007;
  assign n27009 = n7177 & n27008;
  assign n27010 = n8261 & n27009;
  assign n27011 = ~n6784 & n27010;
  assign n27012 = ~n7158 & n27011;
  assign n27013 = ~n8250 & n27012;
  assign n27014 = ~n10642 & n27013;
  assign n27015 = ~n10416 & n27014;
  assign n27016 = ~n9414 & n27015;
  assign n27017 = ~n10641 & n27016;
  assign n27018 = n10640 & n27017;
  assign n27019 = n10638 & n27018;
  assign n27020 = n10666 & n27019;
  assign n27021 = n4955 & n18504;
  assign n27022 = n7909 & n27021;
  assign n27023 = ~n2242 & n27022;
  assign n27024 = ~n3095 & n27023;
  assign n27025 = ~n3997 & n27024;
  assign n27026 = ~n4003 & n27025;
  assign n27027 = ~n4837 & n27026;
  assign n27028 = ~n5822 & n27027;
  assign n27029 = ~n6820 & n27028;
  assign n27030 = ~n7785 & n27029;
  assign n27031 = ~n9027 & n27030;
  assign n27032 = ~n10342 & n27031;
  assign n27033 = ~n10341 & n27032;
  assign n27034 = ~n10245 & n27033;
  assign n27035 = ~n10340 & n27034;
  assign n27036 = n10339 & n27035;
  assign n27037 = n10334 & n27036;
  assign n27038 = n10372 & n27037;
  assign n27039 = ~n27020 & ~n27038;
  assign n27040 = n27006 & n27039;
  assign n27041 = n26981 & n27040;
  assign po105 = ~n26936 | ~n27041;
  assign n27043 = n8363 & n25227;
  assign n27044 = ~n7869 & n27043;
  assign n27045 = ~n8346 & n27044;
  assign n27046 = ~n10714 & n27045;
  assign n27047 = ~n10416 & n27046;
  assign n27048 = ~n9485 & n27047;
  assign n27049 = ~n10713 & n27048;
  assign n27050 = n10640 & n27049;
  assign n27051 = n10712 & n27050;
  assign n27052 = n10740 & n27051;
  assign n27053 = pi105 & ~n4707;
  assign n27054 = n5083 & n27053;
  assign n27055 = n8096 & n27054;
  assign n27056 = n9263 & n27055;
  assign n27057 = ~n4817 & n27056;
  assign n27058 = ~n4902 & n27057;
  assign n27059 = ~n6001 & n27058;
  assign n27060 = ~n7014 & n27059;
  assign n27061 = ~n8114 & n27060;
  assign n27062 = ~n10496 & n27061;
  assign n27063 = ~n10416 & n27062;
  assign n27064 = ~n9276 & n27063;
  assign n27065 = ~n10495 & n27064;
  assign n27066 = n10494 & n27065;
  assign n27067 = n10490 & n27066;
  assign n27068 = n10522 & n27067;
  assign n27069 = ~n27052 & ~n27068;
  assign n27070 = n11378 & n25254;
  assign n27071 = n9942 & n27070;
  assign n27072 = ~n8834 & n27071;
  assign n27073 = ~n11273 & n27072;
  assign n27074 = ~n10416 & n27073;
  assign n27075 = ~n10002 & n27074;
  assign n27076 = ~n10780 & n27075;
  assign n27077 = n10640 & n27076;
  assign n27078 = n11272 & n27077;
  assign n27079 = n11296 & n27078;
  assign n27080 = pi193 & ~n11324;
  assign n27081 = ~n10416 & n27080;
  assign n27082 = ~n10074 & n27081;
  assign n27083 = ~n10780 & n27082;
  assign n27084 = n10640 & n27083;
  assign n27085 = n11323 & n27084;
  assign n27086 = n11342 & n27085;
  assign n27087 = ~n27079 & ~n27086;
  assign n27088 = n27069 & n27087;
  assign n27089 = ~n9215 & n25183;
  assign n27090 = ~n10416 & n27089;
  assign n27091 = ~n10451 & n27090;
  assign n27092 = n10459 & n27091;
  assign n27093 = ~n9160 & n25154;
  assign n27094 = ~n10394 & n27093;
  assign n27095 = n10399 & n27094;
  assign n27096 = pi201 & ~n501;
  assign n27097 = n11440 & n27096;
  assign n27098 = n11446 & n27097;
  assign n27099 = n11437 & n27098;
  assign n27100 = ~n1172 & n27099;
  assign n27101 = ~n996 & n27100;
  assign n27102 = ~n2306 & n27101;
  assign n27103 = ~n500 & n27102;
  assign n27104 = n11004 & n27103;
  assign n27105 = n26550 & n27104;
  assign n27106 = n10980 & n27105;
  assign n27107 = n10971 & n27106;
  assign n27108 = n11172 & n27107;
  assign n27109 = ~n7236 & n27108;
  assign n27110 = ~n6137 & n27109;
  assign n27111 = n6193 & n27110;
  assign n27112 = n6134 & n27111;
  assign n27113 = ~n8867 & n27112;
  assign n27114 = ~n7235 & n27113;
  assign n27115 = n7296 & n27114;
  assign n27116 = n7231 & n27115;
  assign n27117 = ~n10027 & n27116;
  assign n27118 = ~n8866 & n27117;
  assign n27119 = n8898 & n27118;
  assign n27120 = n8863 & n27119;
  assign n27121 = ~n10026 & n27120;
  assign n27122 = n10072 & n27121;
  assign n27123 = n10021 & n27122;
  assign n27124 = pi209 & ~n501;
  assign n27125 = n26571 & n27124;
  assign n27126 = n26575 & n27125;
  assign n27127 = n11404 & n27126;
  assign n27128 = ~n1172 & n27127;
  assign n27129 = ~n996 & n27128;
  assign n27130 = ~n2306 & n27129;
  assign n27131 = ~n500 & n27130;
  assign n27132 = n10855 & n27131;
  assign n27133 = n26584 & n27132;
  assign n27134 = n10831 & n27133;
  assign n27135 = n10823 & n27134;
  assign n27136 = ~n7236 & n27135;
  assign n27137 = ~n6137 & n27136;
  assign n27138 = n6193 & n27137;
  assign n27139 = n6134 & n27138;
  assign n27140 = ~n8867 & n27139;
  assign n27141 = ~n7235 & n27140;
  assign n27142 = n7296 & n27141;
  assign n27143 = n7231 & n27142;
  assign n27144 = ~n10027 & n27143;
  assign n27145 = ~n8866 & n27144;
  assign n27146 = n8898 & n27145;
  assign n27147 = n8863 & n27146;
  assign n27148 = ~n10788 & n27147;
  assign n27149 = ~n10026 & n27148;
  assign n27150 = n10072 & n27149;
  assign n27151 = n10021 & n27150;
  assign n27152 = ~n27123 & ~n27151;
  assign n27153 = ~n27095 & n27152;
  assign n27154 = ~n27092 & n27153;
  assign n27155 = ~n9307 & n25149;
  assign n27156 = ~n10416 & n27155;
  assign n27157 = ~n10452 & n27156;
  assign n27158 = n10552 & n27157;
  assign n27159 = n10546 & n27158;
  assign n27160 = ~n9381 & n25187;
  assign n27161 = ~n10416 & n27160;
  assign n27162 = n10564 & n27161;
  assign n27163 = n10627 & n27162;
  assign n27164 = n10621 & n27163;
  assign n27165 = ~n27159 & ~n27164;
  assign n27166 = n27154 & n27165;
  assign n27167 = pi185 & ~n9687;
  assign n27168 = ~n9913 & n27167;
  assign n27169 = n11365 & n27168;
  assign n27170 = n9856 & n27169;
  assign n27171 = ~n9929 & n27170;
  assign n27172 = ~n10416 & n27171;
  assign n27173 = ~n10622 & n27172;
  assign n27174 = n10564 & n27173;
  assign n27175 = n11226 & n27174;
  assign n27176 = n11218 & n27175;
  assign n27177 = n11265 & n27176;
  assign n27178 = n10602 & n21027;
  assign n27179 = ~n5808 & n27178;
  assign n27180 = ~n6056 & n27179;
  assign n27181 = ~n7073 & n27180;
  assign n27182 = ~n8179 & n27181;
  assign n27183 = ~n10568 & n27182;
  assign n27184 = ~n10416 & n27183;
  assign n27185 = ~n9344 & n27184;
  assign n27186 = ~n10567 & n27185;
  assign n27187 = n10566 & n27186;
  assign n27188 = n10563 & n27187;
  assign n27189 = n10593 & n27188;
  assign n27190 = ~n27177 & ~n27189;
  assign n27191 = n27166 & n27190;
  assign n27192 = n27088 & n27191;
  assign n27193 = pi177 & ~n8900;
  assign n27194 = ~n10416 & n27193;
  assign n27195 = ~n9533 & n27194;
  assign n27196 = ~n10764 & n27195;
  assign n27197 = n10770 & n27196;
  assign n27198 = n10640 & n27197;
  assign n27199 = n10786 & n27198;
  assign n27200 = ~n8397 & n25127;
  assign n27201 = ~n10416 & n27200;
  assign n27202 = ~n10094 & n27201;
  assign n27203 = ~n10713 & n27202;
  assign n27204 = n10640 & n27203;
  assign n27205 = n11312 & n27204;
  assign n27206 = n11305 & n27205;
  assign n27207 = ~n27199 & ~n27206;
  assign n27208 = ~n8291 & n25244;
  assign n27209 = ~n10416 & n27208;
  assign n27210 = ~n9453 & n27209;
  assign n27211 = ~n10696 & n27210;
  assign n27212 = n10702 & n27211;
  assign n27213 = n10640 & n27212;
  assign n27214 = n10695 & n27213;
  assign n27215 = pi041 & ~n1208;
  assign n27216 = n4920 & n27215;
  assign n27217 = n4931 & n27216;
  assign n27218 = n4928 & n27217;
  assign n27219 = ~n1372 & n27218;
  assign n27220 = ~n2243 & n27219;
  assign n27221 = ~n3104 & n27220;
  assign n27222 = ~n3971 & n27221;
  assign n27223 = ~n4003 & n27222;
  assign n27224 = ~n4872 & n27223;
  assign n27225 = ~n5801 & n27224;
  assign n27226 = ~n6739 & n27225;
  assign n27227 = ~n7807 & n27226;
  assign n27228 = ~n8989 & n27227;
  assign n27229 = ~n10293 & n27228;
  assign n27230 = ~n10292 & n27229;
  assign n27231 = ~n10273 & n27230;
  assign n27232 = ~n10291 & n27231;
  assign n27233 = n10290 & n27232;
  assign n27234 = n10285 & n27233;
  assign n27235 = n10326 & n27234;
  assign n27236 = ~n27214 & ~n27235;
  assign n27237 = n27207 & n27236;
  assign n27238 = pi137 & ~n6313;
  assign n27239 = n7169 & n27238;
  assign n27240 = n7177 & n27239;
  assign n27241 = n8261 & n27240;
  assign n27242 = ~n6784 & n27241;
  assign n27243 = ~n7158 & n27242;
  assign n27244 = ~n8250 & n27243;
  assign n27245 = ~n10642 & n27244;
  assign n27246 = ~n10416 & n27245;
  assign n27247 = ~n9414 & n27246;
  assign n27248 = ~n10641 & n27247;
  assign n27249 = n10640 & n27248;
  assign n27250 = n10638 & n27249;
  assign n27251 = n10666 & n27250;
  assign n27252 = n10376 & n25206;
  assign n27253 = n9115 & n27252;
  assign n27254 = ~n3066 & n27253;
  assign n27255 = ~n3983 & n27254;
  assign n27256 = ~n4003 & n27255;
  assign n27257 = ~n4024 & n27256;
  assign n27258 = ~n4999 & n27257;
  assign n27259 = ~n5827 & n27258;
  assign n27260 = ~n6893 & n27259;
  assign n27261 = ~n7890 & n27260;
  assign n27262 = ~n10206 & n27261;
  assign n27263 = ~n10205 & n27262;
  assign n27264 = ~n9131 & n27263;
  assign n27265 = ~n10204 & n27264;
  assign n27266 = n10203 & n27265;
  assign n27267 = n10198 & n27266;
  assign n27268 = n10277 & n27267;
  assign n27269 = ~n27251 & ~n27268;
  assign n27270 = pi089 & ~n3710;
  assign n27271 = n4096 & n27270;
  assign n27272 = n4104 & n27271;
  assign n27273 = n8056 & n27272;
  assign n27274 = ~n3940 & n27273;
  assign n27275 = ~n4001 & n27274;
  assign n27276 = ~n5043 & n27275;
  assign n27277 = ~n5943 & n27276;
  assign n27278 = ~n6951 & n27277;
  assign n27279 = ~n8037 & n27278;
  assign n27280 = ~n10417 & n27279;
  assign n27281 = ~n10416 & n27280;
  assign n27282 = ~n9200 & n27281;
  assign n27283 = ~n10415 & n27282;
  assign n27284 = n10414 & n27283;
  assign n27285 = n10409 & n27284;
  assign n27286 = n10444 & n27285;
  assign n27287 = n4955 & n18542;
  assign n27288 = n7909 & n27287;
  assign n27289 = ~n2242 & n27288;
  assign n27290 = ~n3095 & n27289;
  assign n27291 = ~n3997 & n27290;
  assign n27292 = ~n4003 & n27291;
  assign n27293 = ~n4837 & n27292;
  assign n27294 = ~n5822 & n27293;
  assign n27295 = ~n6820 & n27294;
  assign n27296 = ~n7785 & n27295;
  assign n27297 = ~n9027 & n27296;
  assign n27298 = ~n10342 & n27297;
  assign n27299 = ~n10341 & n27298;
  assign n27300 = ~n10245 & n27299;
  assign n27301 = ~n10340 & n27300;
  assign n27302 = n10339 & n27301;
  assign n27303 = n10334 & n27302;
  assign n27304 = n10372 & n27303;
  assign n27305 = ~n27286 & ~n27304;
  assign n27306 = n27269 & n27305;
  assign n27307 = n27237 & n27306;
  assign po106 = ~n27192 | ~n27307;
  assign n27309 = n8363 & n25458;
  assign n27310 = ~n7869 & n27309;
  assign n27311 = ~n8346 & n27310;
  assign n27312 = ~n10714 & n27311;
  assign n27313 = ~n10416 & n27312;
  assign n27314 = ~n9485 & n27313;
  assign n27315 = ~n10713 & n27314;
  assign n27316 = n10640 & n27315;
  assign n27317 = n10712 & n27316;
  assign n27318 = n10740 & n27317;
  assign n27319 = n10376 & n25413;
  assign n27320 = n9115 & n27319;
  assign n27321 = ~n3066 & n27320;
  assign n27322 = ~n3983 & n27321;
  assign n27323 = ~n4003 & n27322;
  assign n27324 = ~n4024 & n27323;
  assign n27325 = ~n4999 & n27324;
  assign n27326 = ~n5827 & n27325;
  assign n27327 = ~n6893 & n27326;
  assign n27328 = ~n7890 & n27327;
  assign n27329 = ~n10206 & n27328;
  assign n27330 = ~n10205 & n27329;
  assign n27331 = ~n9131 & n27330;
  assign n27332 = ~n10204 & n27331;
  assign n27333 = n10203 & n27332;
  assign n27334 = n10198 & n27333;
  assign n27335 = n10277 & n27334;
  assign n27336 = ~n27318 & ~n27335;
  assign n27337 = ~n8397 & n25315;
  assign n27338 = ~n10416 & n27337;
  assign n27339 = ~n10094 & n27338;
  assign n27340 = ~n10713 & n27339;
  assign n27341 = n10640 & n27340;
  assign n27342 = n11312 & n27341;
  assign n27343 = n11305 & n27342;
  assign n27344 = pi186 & ~n9687;
  assign n27345 = ~n9913 & n27344;
  assign n27346 = n11365 & n27345;
  assign n27347 = n9856 & n27346;
  assign n27348 = ~n9929 & n27347;
  assign n27349 = ~n10416 & n27348;
  assign n27350 = ~n10622 & n27349;
  assign n27351 = n10564 & n27350;
  assign n27352 = n11226 & n27351;
  assign n27353 = n11218 & n27352;
  assign n27354 = n11265 & n27353;
  assign n27355 = ~n27343 & ~n27354;
  assign n27356 = n27336 & n27355;
  assign n27357 = ~n9215 & n25390;
  assign n27358 = ~n10416 & n27357;
  assign n27359 = ~n10451 & n27358;
  assign n27360 = n10459 & n27359;
  assign n27361 = ~n9160 & n25361;
  assign n27362 = ~n10394 & n27361;
  assign n27363 = n10399 & n27362;
  assign n27364 = pi202 & ~n501;
  assign n27365 = n11440 & n27364;
  assign n27366 = n11446 & n27365;
  assign n27367 = n11437 & n27366;
  assign n27368 = ~n1172 & n27367;
  assign n27369 = ~n996 & n27368;
  assign n27370 = ~n2306 & n27369;
  assign n27371 = ~n500 & n27370;
  assign n27372 = n11004 & n27371;
  assign n27373 = n26550 & n27372;
  assign n27374 = n10980 & n27373;
  assign n27375 = n10971 & n27374;
  assign n27376 = n11172 & n27375;
  assign n27377 = ~n7236 & n27376;
  assign n27378 = ~n6137 & n27377;
  assign n27379 = n6193 & n27378;
  assign n27380 = n6134 & n27379;
  assign n27381 = ~n8867 & n27380;
  assign n27382 = ~n7235 & n27381;
  assign n27383 = n7296 & n27382;
  assign n27384 = n7231 & n27383;
  assign n27385 = ~n10027 & n27384;
  assign n27386 = ~n8866 & n27385;
  assign n27387 = n8898 & n27386;
  assign n27388 = n8863 & n27387;
  assign n27389 = ~n10026 & n27388;
  assign n27390 = n10072 & n27389;
  assign n27391 = n10021 & n27390;
  assign n27392 = pi210 & ~n501;
  assign n27393 = n26571 & n27392;
  assign n27394 = n26575 & n27393;
  assign n27395 = n11404 & n27394;
  assign n27396 = ~n1172 & n27395;
  assign n27397 = ~n996 & n27396;
  assign n27398 = ~n2306 & n27397;
  assign n27399 = ~n500 & n27398;
  assign n27400 = n10855 & n27399;
  assign n27401 = n26584 & n27400;
  assign n27402 = n10831 & n27401;
  assign n27403 = n10823 & n27402;
  assign n27404 = ~n7236 & n27403;
  assign n27405 = ~n6137 & n27404;
  assign n27406 = n6193 & n27405;
  assign n27407 = n6134 & n27406;
  assign n27408 = ~n8867 & n27407;
  assign n27409 = ~n7235 & n27408;
  assign n27410 = n7296 & n27409;
  assign n27411 = n7231 & n27410;
  assign n27412 = ~n10027 & n27411;
  assign n27413 = ~n8866 & n27412;
  assign n27414 = n8898 & n27413;
  assign n27415 = n8863 & n27414;
  assign n27416 = ~n10788 & n27415;
  assign n27417 = ~n10026 & n27416;
  assign n27418 = n10072 & n27417;
  assign n27419 = n10021 & n27418;
  assign n27420 = ~n27391 & ~n27419;
  assign n27421 = ~n27363 & n27420;
  assign n27422 = ~n27360 & n27421;
  assign n27423 = ~n9307 & n25356;
  assign n27424 = ~n10416 & n27423;
  assign n27425 = ~n10452 & n27424;
  assign n27426 = n10552 & n27425;
  assign n27427 = n10546 & n27426;
  assign n27428 = ~n9381 & n25394;
  assign n27429 = ~n10416 & n27428;
  assign n27430 = n10564 & n27429;
  assign n27431 = n10627 & n27430;
  assign n27432 = n10621 & n27431;
  assign n27433 = ~n27427 & ~n27432;
  assign n27434 = n27422 & n27433;
  assign n27435 = pi138 & ~n6313;
  assign n27436 = n7169 & n27435;
  assign n27437 = n7177 & n27436;
  assign n27438 = n8261 & n27437;
  assign n27439 = ~n6784 & n27438;
  assign n27440 = ~n7158 & n27439;
  assign n27441 = ~n8250 & n27440;
  assign n27442 = ~n10642 & n27441;
  assign n27443 = ~n10416 & n27442;
  assign n27444 = ~n9414 & n27443;
  assign n27445 = ~n10641 & n27444;
  assign n27446 = n10640 & n27445;
  assign n27447 = n10638 & n27446;
  assign n27448 = n10666 & n27447;
  assign n27449 = n4955 & n18580;
  assign n27450 = n7909 & n27449;
  assign n27451 = ~n2242 & n27450;
  assign n27452 = ~n3095 & n27451;
  assign n27453 = ~n3997 & n27452;
  assign n27454 = ~n4003 & n27453;
  assign n27455 = ~n4837 & n27454;
  assign n27456 = ~n5822 & n27455;
  assign n27457 = ~n6820 & n27456;
  assign n27458 = ~n7785 & n27457;
  assign n27459 = ~n9027 & n27458;
  assign n27460 = ~n10342 & n27459;
  assign n27461 = ~n10341 & n27460;
  assign n27462 = ~n10245 & n27461;
  assign n27463 = ~n10340 & n27462;
  assign n27464 = n10339 & n27463;
  assign n27465 = n10334 & n27464;
  assign n27466 = n10372 & n27465;
  assign n27467 = ~n27448 & ~n27466;
  assign n27468 = n27434 & n27467;
  assign n27469 = n27356 & n27468;
  assign n27470 = ~n8291 & n25347;
  assign n27471 = ~n10416 & n27470;
  assign n27472 = ~n9453 & n27471;
  assign n27473 = ~n10696 & n27472;
  assign n27474 = n10702 & n27473;
  assign n27475 = n10640 & n27474;
  assign n27476 = n10695 & n27475;
  assign n27477 = pi042 & ~n1208;
  assign n27478 = n4920 & n27477;
  assign n27479 = n4931 & n27478;
  assign n27480 = n4928 & n27479;
  assign n27481 = ~n1372 & n27480;
  assign n27482 = ~n2243 & n27481;
  assign n27483 = ~n3104 & n27482;
  assign n27484 = ~n3971 & n27483;
  assign n27485 = ~n4003 & n27484;
  assign n27486 = ~n4872 & n27485;
  assign n27487 = ~n5801 & n27486;
  assign n27488 = ~n6739 & n27487;
  assign n27489 = ~n7807 & n27488;
  assign n27490 = ~n8989 & n27489;
  assign n27491 = ~n10293 & n27490;
  assign n27492 = ~n10292 & n27491;
  assign n27493 = ~n10273 & n27492;
  assign n27494 = ~n10291 & n27493;
  assign n27495 = n10290 & n27494;
  assign n27496 = n10285 & n27495;
  assign n27497 = n10326 & n27496;
  assign n27498 = ~n27476 & ~n27497;
  assign n27499 = pi178 & ~n8900;
  assign n27500 = ~n10416 & n27499;
  assign n27501 = ~n9533 & n27500;
  assign n27502 = ~n10764 & n27501;
  assign n27503 = n10770 & n27502;
  assign n27504 = n10640 & n27503;
  assign n27505 = n10786 & n27504;
  assign n27506 = pi090 & ~n3710;
  assign n27507 = n4096 & n27506;
  assign n27508 = n4104 & n27507;
  assign n27509 = n8056 & n27508;
  assign n27510 = ~n3940 & n27509;
  assign n27511 = ~n4001 & n27510;
  assign n27512 = ~n5043 & n27511;
  assign n27513 = ~n5943 & n27512;
  assign n27514 = ~n6951 & n27513;
  assign n27515 = ~n8037 & n27514;
  assign n27516 = ~n10417 & n27515;
  assign n27517 = ~n10416 & n27516;
  assign n27518 = ~n9200 & n27517;
  assign n27519 = ~n10415 & n27518;
  assign n27520 = n10414 & n27519;
  assign n27521 = n10409 & n27520;
  assign n27522 = n10444 & n27521;
  assign n27523 = ~n27505 & ~n27522;
  assign n27524 = n27498 & n27523;
  assign n27525 = n10602 & n21153;
  assign n27526 = ~n5808 & n27525;
  assign n27527 = ~n6056 & n27526;
  assign n27528 = ~n7073 & n27527;
  assign n27529 = ~n8179 & n27528;
  assign n27530 = ~n10568 & n27529;
  assign n27531 = ~n10416 & n27530;
  assign n27532 = ~n9344 & n27531;
  assign n27533 = ~n10567 & n27532;
  assign n27534 = n10566 & n27533;
  assign n27535 = n10563 & n27534;
  assign n27536 = n10593 & n27535;
  assign n27537 = pi106 & ~n4707;
  assign n27538 = n5083 & n27537;
  assign n27539 = n8096 & n27538;
  assign n27540 = n9263 & n27539;
  assign n27541 = ~n4817 & n27540;
  assign n27542 = ~n4902 & n27541;
  assign n27543 = ~n6001 & n27542;
  assign n27544 = ~n7014 & n27543;
  assign n27545 = ~n8114 & n27544;
  assign n27546 = ~n10496 & n27545;
  assign n27547 = ~n10416 & n27546;
  assign n27548 = ~n9276 & n27547;
  assign n27549 = ~n10495 & n27548;
  assign n27550 = n10494 & n27549;
  assign n27551 = n10490 & n27550;
  assign n27552 = n10522 & n27551;
  assign n27553 = ~n27536 & ~n27552;
  assign n27554 = n11378 & n25514;
  assign n27555 = n9942 & n27554;
  assign n27556 = ~n8834 & n27555;
  assign n27557 = ~n11273 & n27556;
  assign n27558 = ~n10416 & n27557;
  assign n27559 = ~n10002 & n27558;
  assign n27560 = ~n10780 & n27559;
  assign n27561 = n10640 & n27560;
  assign n27562 = n11272 & n27561;
  assign n27563 = n11296 & n27562;
  assign n27564 = pi194 & ~n11324;
  assign n27565 = ~n10416 & n27564;
  assign n27566 = ~n10074 & n27565;
  assign n27567 = ~n10780 & n27566;
  assign n27568 = n10640 & n27567;
  assign n27569 = n11323 & n27568;
  assign n27570 = n11342 & n27569;
  assign n27571 = ~n27563 & ~n27570;
  assign n27572 = n27553 & n27571;
  assign n27573 = n27524 & n27572;
  assign po107 = ~n27469 | ~n27573;
  assign n27575 = n4955 & n18618;
  assign n27576 = n7909 & n27575;
  assign n27577 = ~n2242 & n27576;
  assign n27578 = ~n3095 & n27577;
  assign n27579 = ~n3997 & n27578;
  assign n27580 = ~n4003 & n27579;
  assign n27581 = ~n4837 & n27580;
  assign n27582 = ~n5822 & n27581;
  assign n27583 = ~n6820 & n27582;
  assign n27584 = ~n7785 & n27583;
  assign n27585 = ~n9027 & n27584;
  assign n27586 = ~n10342 & n27585;
  assign n27587 = ~n10341 & n27586;
  assign n27588 = ~n10245 & n27587;
  assign n27589 = ~n10340 & n27588;
  assign n27590 = n10339 & n27589;
  assign n27591 = n10334 & n27590;
  assign n27592 = n10372 & n27591;
  assign n27593 = pi179 & ~n8900;
  assign n27594 = ~n10416 & n27593;
  assign n27595 = ~n9533 & n27594;
  assign n27596 = ~n10764 & n27595;
  assign n27597 = n10770 & n27596;
  assign n27598 = n10640 & n27597;
  assign n27599 = n10786 & n27598;
  assign n27600 = ~n27592 & ~n27599;
  assign n27601 = ~n8397 & n25745;
  assign n27602 = ~n10416 & n27601;
  assign n27603 = ~n10094 & n27602;
  assign n27604 = ~n10713 & n27603;
  assign n27605 = n10640 & n27604;
  assign n27606 = n11312 & n27605;
  assign n27607 = n11305 & n27606;
  assign n27608 = pi187 & ~n9687;
  assign n27609 = ~n9913 & n27608;
  assign n27610 = n11365 & n27609;
  assign n27611 = n9856 & n27610;
  assign n27612 = ~n9929 & n27611;
  assign n27613 = ~n10416 & n27612;
  assign n27614 = ~n10622 & n27613;
  assign n27615 = n10564 & n27614;
  assign n27616 = n11226 & n27615;
  assign n27617 = n11218 & n27616;
  assign n27618 = n11265 & n27617;
  assign n27619 = ~n27607 & ~n27618;
  assign n27620 = n27600 & n27619;
  assign n27621 = ~n9215 & n25647;
  assign n27622 = ~n10416 & n27621;
  assign n27623 = ~n10451 & n27622;
  assign n27624 = n10459 & n27623;
  assign n27625 = ~n9160 & n25618;
  assign n27626 = ~n10394 & n27625;
  assign n27627 = n10399 & n27626;
  assign n27628 = pi203 & ~n501;
  assign n27629 = n11440 & n27628;
  assign n27630 = n11446 & n27629;
  assign n27631 = n11437 & n27630;
  assign n27632 = ~n1172 & n27631;
  assign n27633 = ~n996 & n27632;
  assign n27634 = ~n2306 & n27633;
  assign n27635 = ~n500 & n27634;
  assign n27636 = n11004 & n27635;
  assign n27637 = n26550 & n27636;
  assign n27638 = n10980 & n27637;
  assign n27639 = n10971 & n27638;
  assign n27640 = n11172 & n27639;
  assign n27641 = ~n7236 & n27640;
  assign n27642 = ~n6137 & n27641;
  assign n27643 = n6193 & n27642;
  assign n27644 = n6134 & n27643;
  assign n27645 = ~n8867 & n27644;
  assign n27646 = ~n7235 & n27645;
  assign n27647 = n7296 & n27646;
  assign n27648 = n7231 & n27647;
  assign n27649 = ~n10027 & n27648;
  assign n27650 = ~n8866 & n27649;
  assign n27651 = n8898 & n27650;
  assign n27652 = n8863 & n27651;
  assign n27653 = ~n10026 & n27652;
  assign n27654 = n10072 & n27653;
  assign n27655 = n10021 & n27654;
  assign n27656 = pi211 & ~n501;
  assign n27657 = n26571 & n27656;
  assign n27658 = n26575 & n27657;
  assign n27659 = n11404 & n27658;
  assign n27660 = ~n1172 & n27659;
  assign n27661 = ~n996 & n27660;
  assign n27662 = ~n2306 & n27661;
  assign n27663 = ~n500 & n27662;
  assign n27664 = n10855 & n27663;
  assign n27665 = n26584 & n27664;
  assign n27666 = n10831 & n27665;
  assign n27667 = n10823 & n27666;
  assign n27668 = ~n7236 & n27667;
  assign n27669 = ~n6137 & n27668;
  assign n27670 = n6193 & n27669;
  assign n27671 = n6134 & n27670;
  assign n27672 = ~n8867 & n27671;
  assign n27673 = ~n7235 & n27672;
  assign n27674 = n7296 & n27673;
  assign n27675 = n7231 & n27674;
  assign n27676 = ~n10027 & n27675;
  assign n27677 = ~n8866 & n27676;
  assign n27678 = n8898 & n27677;
  assign n27679 = n8863 & n27678;
  assign n27680 = ~n10788 & n27679;
  assign n27681 = ~n10026 & n27680;
  assign n27682 = n10072 & n27681;
  assign n27683 = n10021 & n27682;
  assign n27684 = ~n27655 & ~n27683;
  assign n27685 = ~n27627 & n27684;
  assign n27686 = ~n27624 & n27685;
  assign n27687 = ~n9307 & n25613;
  assign n27688 = ~n10416 & n27687;
  assign n27689 = ~n10452 & n27688;
  assign n27690 = n10552 & n27689;
  assign n27691 = n10546 & n27690;
  assign n27692 = ~n9381 & n25651;
  assign n27693 = ~n10416 & n27692;
  assign n27694 = n10564 & n27693;
  assign n27695 = n10627 & n27694;
  assign n27696 = n10621 & n27695;
  assign n27697 = ~n27691 & ~n27696;
  assign n27698 = n27686 & n27697;
  assign n27699 = n8363 & n25576;
  assign n27700 = ~n7869 & n27699;
  assign n27701 = ~n8346 & n27700;
  assign n27702 = ~n10714 & n27701;
  assign n27703 = ~n10416 & n27702;
  assign n27704 = ~n9485 & n27703;
  assign n27705 = ~n10713 & n27704;
  assign n27706 = n10640 & n27705;
  assign n27707 = n10712 & n27706;
  assign n27708 = n10740 & n27707;
  assign n27709 = n10602 & n21279;
  assign n27710 = ~n5808 & n27709;
  assign n27711 = ~n6056 & n27710;
  assign n27712 = ~n7073 & n27711;
  assign n27713 = ~n8179 & n27712;
  assign n27714 = ~n10568 & n27713;
  assign n27715 = ~n10416 & n27714;
  assign n27716 = ~n9344 & n27715;
  assign n27717 = ~n10567 & n27716;
  assign n27718 = n10566 & n27717;
  assign n27719 = n10563 & n27718;
  assign n27720 = n10593 & n27719;
  assign n27721 = ~n27708 & ~n27720;
  assign n27722 = n27698 & n27721;
  assign n27723 = n27620 & n27722;
  assign n27724 = ~n8291 & n25701;
  assign n27725 = ~n10416 & n27724;
  assign n27726 = ~n9453 & n27725;
  assign n27727 = ~n10696 & n27726;
  assign n27728 = n10702 & n27727;
  assign n27729 = n10640 & n27728;
  assign n27730 = n10695 & n27729;
  assign n27731 = pi043 & ~n1208;
  assign n27732 = n4920 & n27731;
  assign n27733 = n4931 & n27732;
  assign n27734 = n4928 & n27733;
  assign n27735 = ~n1372 & n27734;
  assign n27736 = ~n2243 & n27735;
  assign n27737 = ~n3104 & n27736;
  assign n27738 = ~n3971 & n27737;
  assign n27739 = ~n4003 & n27738;
  assign n27740 = ~n4872 & n27739;
  assign n27741 = ~n5801 & n27740;
  assign n27742 = ~n6739 & n27741;
  assign n27743 = ~n7807 & n27742;
  assign n27744 = ~n8989 & n27743;
  assign n27745 = ~n10293 & n27744;
  assign n27746 = ~n10292 & n27745;
  assign n27747 = ~n10273 & n27746;
  assign n27748 = ~n10291 & n27747;
  assign n27749 = n10290 & n27748;
  assign n27750 = n10285 & n27749;
  assign n27751 = n10326 & n27750;
  assign n27752 = ~n27730 & ~n27751;
  assign n27753 = n10376 & n25670;
  assign n27754 = n9115 & n27753;
  assign n27755 = ~n3066 & n27754;
  assign n27756 = ~n3983 & n27755;
  assign n27757 = ~n4003 & n27756;
  assign n27758 = ~n4024 & n27757;
  assign n27759 = ~n4999 & n27758;
  assign n27760 = ~n5827 & n27759;
  assign n27761 = ~n6893 & n27760;
  assign n27762 = ~n7890 & n27761;
  assign n27763 = ~n10206 & n27762;
  assign n27764 = ~n10205 & n27763;
  assign n27765 = ~n9131 & n27764;
  assign n27766 = ~n10204 & n27765;
  assign n27767 = n10203 & n27766;
  assign n27768 = n10198 & n27767;
  assign n27769 = n10277 & n27768;
  assign n27770 = pi091 & ~n3710;
  assign n27771 = n4096 & n27770;
  assign n27772 = n4104 & n27771;
  assign n27773 = n8056 & n27772;
  assign n27774 = ~n3940 & n27773;
  assign n27775 = ~n4001 & n27774;
  assign n27776 = ~n5043 & n27775;
  assign n27777 = ~n5943 & n27776;
  assign n27778 = ~n6951 & n27777;
  assign n27779 = ~n8037 & n27778;
  assign n27780 = ~n10417 & n27779;
  assign n27781 = ~n10416 & n27780;
  assign n27782 = ~n9200 & n27781;
  assign n27783 = ~n10415 & n27782;
  assign n27784 = n10414 & n27783;
  assign n27785 = n10409 & n27784;
  assign n27786 = n10444 & n27785;
  assign n27787 = ~n27769 & ~n27786;
  assign n27788 = n27752 & n27787;
  assign n27789 = pi139 & ~n6313;
  assign n27790 = n7169 & n27789;
  assign n27791 = n7177 & n27790;
  assign n27792 = n8261 & n27791;
  assign n27793 = ~n6784 & n27792;
  assign n27794 = ~n7158 & n27793;
  assign n27795 = ~n8250 & n27794;
  assign n27796 = ~n10642 & n27795;
  assign n27797 = ~n10416 & n27796;
  assign n27798 = ~n9414 & n27797;
  assign n27799 = ~n10641 & n27798;
  assign n27800 = n10640 & n27799;
  assign n27801 = n10638 & n27800;
  assign n27802 = n10666 & n27801;
  assign n27803 = pi107 & ~n4707;
  assign n27804 = n5083 & n27803;
  assign n27805 = n8096 & n27804;
  assign n27806 = n9263 & n27805;
  assign n27807 = ~n4817 & n27806;
  assign n27808 = ~n4902 & n27807;
  assign n27809 = ~n6001 & n27808;
  assign n27810 = ~n7014 & n27809;
  assign n27811 = ~n8114 & n27810;
  assign n27812 = ~n10496 & n27811;
  assign n27813 = ~n10416 & n27812;
  assign n27814 = ~n9276 & n27813;
  assign n27815 = ~n10495 & n27814;
  assign n27816 = n10494 & n27815;
  assign n27817 = n10490 & n27816;
  assign n27818 = n10522 & n27817;
  assign n27819 = ~n27802 & ~n27818;
  assign n27820 = n11378 & n25601;
  assign n27821 = n9942 & n27820;
  assign n27822 = ~n8834 & n27821;
  assign n27823 = ~n11273 & n27822;
  assign n27824 = ~n10416 & n27823;
  assign n27825 = ~n10002 & n27824;
  assign n27826 = ~n10780 & n27825;
  assign n27827 = n10640 & n27826;
  assign n27828 = n11272 & n27827;
  assign n27829 = n11296 & n27828;
  assign n27830 = pi195 & ~n11324;
  assign n27831 = ~n10416 & n27830;
  assign n27832 = ~n10074 & n27831;
  assign n27833 = ~n10780 & n27832;
  assign n27834 = n10640 & n27833;
  assign n27835 = n11323 & n27834;
  assign n27836 = n11342 & n27835;
  assign n27837 = ~n27829 & ~n27836;
  assign n27838 = n27819 & n27837;
  assign n27839 = n27788 & n27838;
  assign po108 = ~n27723 | ~n27839;
  assign n27841 = n4955 & n18656;
  assign n27842 = n7909 & n27841;
  assign n27843 = ~n2242 & n27842;
  assign n27844 = ~n3095 & n27843;
  assign n27845 = ~n3997 & n27844;
  assign n27846 = ~n4003 & n27845;
  assign n27847 = ~n4837 & n27846;
  assign n27848 = ~n5822 & n27847;
  assign n27849 = ~n6820 & n27848;
  assign n27850 = ~n7785 & n27849;
  assign n27851 = ~n9027 & n27850;
  assign n27852 = ~n10342 & n27851;
  assign n27853 = ~n10341 & n27852;
  assign n27854 = ~n10245 & n27853;
  assign n27855 = ~n10340 & n27854;
  assign n27856 = n10339 & n27855;
  assign n27857 = n10334 & n27856;
  assign n27858 = n10372 & n27857;
  assign n27859 = pi180 & ~n8900;
  assign n27860 = ~n10416 & n27859;
  assign n27861 = ~n9533 & n27860;
  assign n27862 = ~n10764 & n27861;
  assign n27863 = n10770 & n27862;
  assign n27864 = n10640 & n27863;
  assign n27865 = n10786 & n27864;
  assign n27866 = ~n27858 & ~n27865;
  assign n27867 = ~n8397 & n25978;
  assign n27868 = ~n10416 & n27867;
  assign n27869 = ~n10094 & n27868;
  assign n27870 = ~n10713 & n27869;
  assign n27871 = n10640 & n27870;
  assign n27872 = n11312 & n27871;
  assign n27873 = n11305 & n27872;
  assign n27874 = pi188 & ~n9687;
  assign n27875 = ~n9913 & n27874;
  assign n27876 = n11365 & n27875;
  assign n27877 = n9856 & n27876;
  assign n27878 = ~n9929 & n27877;
  assign n27879 = ~n10416 & n27878;
  assign n27880 = ~n10622 & n27879;
  assign n27881 = n10564 & n27880;
  assign n27882 = n11226 & n27881;
  assign n27883 = n11218 & n27882;
  assign n27884 = n11265 & n27883;
  assign n27885 = ~n27873 & ~n27884;
  assign n27886 = n27866 & n27885;
  assign n27887 = ~n9215 & n25880;
  assign n27888 = ~n10416 & n27887;
  assign n27889 = ~n10451 & n27888;
  assign n27890 = n10459 & n27889;
  assign n27891 = ~n9160 & n25851;
  assign n27892 = ~n10394 & n27891;
  assign n27893 = n10399 & n27892;
  assign n27894 = pi204 & ~n501;
  assign n27895 = n11440 & n27894;
  assign n27896 = n11446 & n27895;
  assign n27897 = n11437 & n27896;
  assign n27898 = ~n1172 & n27897;
  assign n27899 = ~n996 & n27898;
  assign n27900 = ~n2306 & n27899;
  assign n27901 = ~n500 & n27900;
  assign n27902 = n11004 & n27901;
  assign n27903 = n26550 & n27902;
  assign n27904 = n10980 & n27903;
  assign n27905 = n10971 & n27904;
  assign n27906 = n11172 & n27905;
  assign n27907 = ~n7236 & n27906;
  assign n27908 = ~n6137 & n27907;
  assign n27909 = n6193 & n27908;
  assign n27910 = n6134 & n27909;
  assign n27911 = ~n8867 & n27910;
  assign n27912 = ~n7235 & n27911;
  assign n27913 = n7296 & n27912;
  assign n27914 = n7231 & n27913;
  assign n27915 = ~n10027 & n27914;
  assign n27916 = ~n8866 & n27915;
  assign n27917 = n8898 & n27916;
  assign n27918 = n8863 & n27917;
  assign n27919 = ~n10026 & n27918;
  assign n27920 = n10072 & n27919;
  assign n27921 = n10021 & n27920;
  assign n27922 = pi212 & ~n501;
  assign n27923 = n26571 & n27922;
  assign n27924 = n26575 & n27923;
  assign n27925 = n11404 & n27924;
  assign n27926 = ~n1172 & n27925;
  assign n27927 = ~n996 & n27926;
  assign n27928 = ~n2306 & n27927;
  assign n27929 = ~n500 & n27928;
  assign n27930 = n10855 & n27929;
  assign n27931 = n26584 & n27930;
  assign n27932 = n10831 & n27931;
  assign n27933 = n10823 & n27932;
  assign n27934 = ~n7236 & n27933;
  assign n27935 = ~n6137 & n27934;
  assign n27936 = n6193 & n27935;
  assign n27937 = n6134 & n27936;
  assign n27938 = ~n8867 & n27937;
  assign n27939 = ~n7235 & n27938;
  assign n27940 = n7296 & n27939;
  assign n27941 = n7231 & n27940;
  assign n27942 = ~n10027 & n27941;
  assign n27943 = ~n8866 & n27942;
  assign n27944 = n8898 & n27943;
  assign n27945 = n8863 & n27944;
  assign n27946 = ~n10788 & n27945;
  assign n27947 = ~n10026 & n27946;
  assign n27948 = n10072 & n27947;
  assign n27949 = n10021 & n27948;
  assign n27950 = ~n27921 & ~n27949;
  assign n27951 = ~n27893 & n27950;
  assign n27952 = ~n27890 & n27951;
  assign n27953 = ~n9307 & n25846;
  assign n27954 = ~n10416 & n27953;
  assign n27955 = ~n10452 & n27954;
  assign n27956 = n10552 & n27955;
  assign n27957 = n10546 & n27956;
  assign n27958 = ~n9381 & n25884;
  assign n27959 = ~n10416 & n27958;
  assign n27960 = n10564 & n27959;
  assign n27961 = n10627 & n27960;
  assign n27962 = n10621 & n27961;
  assign n27963 = ~n27957 & ~n27962;
  assign n27964 = n27952 & n27963;
  assign n27965 = n8363 & n25809;
  assign n27966 = ~n7869 & n27965;
  assign n27967 = ~n8346 & n27966;
  assign n27968 = ~n10714 & n27967;
  assign n27969 = ~n10416 & n27968;
  assign n27970 = ~n9485 & n27969;
  assign n27971 = ~n10713 & n27970;
  assign n27972 = n10640 & n27971;
  assign n27973 = n10712 & n27972;
  assign n27974 = n10740 & n27973;
  assign n27975 = n10602 & n21405;
  assign n27976 = ~n5808 & n27975;
  assign n27977 = ~n6056 & n27976;
  assign n27978 = ~n7073 & n27977;
  assign n27979 = ~n8179 & n27978;
  assign n27980 = ~n10568 & n27979;
  assign n27981 = ~n10416 & n27980;
  assign n27982 = ~n9344 & n27981;
  assign n27983 = ~n10567 & n27982;
  assign n27984 = n10566 & n27983;
  assign n27985 = n10563 & n27984;
  assign n27986 = n10593 & n27985;
  assign n27987 = ~n27974 & ~n27986;
  assign n27988 = n27964 & n27987;
  assign n27989 = n27886 & n27988;
  assign n27990 = ~n8291 & n25934;
  assign n27991 = ~n10416 & n27990;
  assign n27992 = ~n9453 & n27991;
  assign n27993 = ~n10696 & n27992;
  assign n27994 = n10702 & n27993;
  assign n27995 = n10640 & n27994;
  assign n27996 = n10695 & n27995;
  assign n27997 = pi044 & ~n1208;
  assign n27998 = n4920 & n27997;
  assign n27999 = n4931 & n27998;
  assign n28000 = n4928 & n27999;
  assign n28001 = ~n1372 & n28000;
  assign n28002 = ~n2243 & n28001;
  assign n28003 = ~n3104 & n28002;
  assign n28004 = ~n3971 & n28003;
  assign n28005 = ~n4003 & n28004;
  assign n28006 = ~n4872 & n28005;
  assign n28007 = ~n5801 & n28006;
  assign n28008 = ~n6739 & n28007;
  assign n28009 = ~n7807 & n28008;
  assign n28010 = ~n8989 & n28009;
  assign n28011 = ~n10293 & n28010;
  assign n28012 = ~n10292 & n28011;
  assign n28013 = ~n10273 & n28012;
  assign n28014 = ~n10291 & n28013;
  assign n28015 = n10290 & n28014;
  assign n28016 = n10285 & n28015;
  assign n28017 = n10326 & n28016;
  assign n28018 = ~n27996 & ~n28017;
  assign n28019 = n10376 & n25903;
  assign n28020 = n9115 & n28019;
  assign n28021 = ~n3066 & n28020;
  assign n28022 = ~n3983 & n28021;
  assign n28023 = ~n4003 & n28022;
  assign n28024 = ~n4024 & n28023;
  assign n28025 = ~n4999 & n28024;
  assign n28026 = ~n5827 & n28025;
  assign n28027 = ~n6893 & n28026;
  assign n28028 = ~n7890 & n28027;
  assign n28029 = ~n10206 & n28028;
  assign n28030 = ~n10205 & n28029;
  assign n28031 = ~n9131 & n28030;
  assign n28032 = ~n10204 & n28031;
  assign n28033 = n10203 & n28032;
  assign n28034 = n10198 & n28033;
  assign n28035 = n10277 & n28034;
  assign n28036 = pi092 & ~n3710;
  assign n28037 = n4096 & n28036;
  assign n28038 = n4104 & n28037;
  assign n28039 = n8056 & n28038;
  assign n28040 = ~n3940 & n28039;
  assign n28041 = ~n4001 & n28040;
  assign n28042 = ~n5043 & n28041;
  assign n28043 = ~n5943 & n28042;
  assign n28044 = ~n6951 & n28043;
  assign n28045 = ~n8037 & n28044;
  assign n28046 = ~n10417 & n28045;
  assign n28047 = ~n10416 & n28046;
  assign n28048 = ~n9200 & n28047;
  assign n28049 = ~n10415 & n28048;
  assign n28050 = n10414 & n28049;
  assign n28051 = n10409 & n28050;
  assign n28052 = n10444 & n28051;
  assign n28053 = ~n28035 & ~n28052;
  assign n28054 = n28018 & n28053;
  assign n28055 = pi140 & ~n6313;
  assign n28056 = n7169 & n28055;
  assign n28057 = n7177 & n28056;
  assign n28058 = n8261 & n28057;
  assign n28059 = ~n6784 & n28058;
  assign n28060 = ~n7158 & n28059;
  assign n28061 = ~n8250 & n28060;
  assign n28062 = ~n10642 & n28061;
  assign n28063 = ~n10416 & n28062;
  assign n28064 = ~n9414 & n28063;
  assign n28065 = ~n10641 & n28064;
  assign n28066 = n10640 & n28065;
  assign n28067 = n10638 & n28066;
  assign n28068 = n10666 & n28067;
  assign n28069 = pi108 & ~n4707;
  assign n28070 = n5083 & n28069;
  assign n28071 = n8096 & n28070;
  assign n28072 = n9263 & n28071;
  assign n28073 = ~n4817 & n28072;
  assign n28074 = ~n4902 & n28073;
  assign n28075 = ~n6001 & n28074;
  assign n28076 = ~n7014 & n28075;
  assign n28077 = ~n8114 & n28076;
  assign n28078 = ~n10496 & n28077;
  assign n28079 = ~n10416 & n28078;
  assign n28080 = ~n9276 & n28079;
  assign n28081 = ~n10495 & n28080;
  assign n28082 = n10494 & n28081;
  assign n28083 = n10490 & n28082;
  assign n28084 = n10522 & n28083;
  assign n28085 = ~n28068 & ~n28084;
  assign n28086 = n11378 & n25834;
  assign n28087 = n9942 & n28086;
  assign n28088 = ~n8834 & n28087;
  assign n28089 = ~n11273 & n28088;
  assign n28090 = ~n10416 & n28089;
  assign n28091 = ~n10002 & n28090;
  assign n28092 = ~n10780 & n28091;
  assign n28093 = n10640 & n28092;
  assign n28094 = n11272 & n28093;
  assign n28095 = n11296 & n28094;
  assign n28096 = pi196 & ~n11324;
  assign n28097 = ~n10416 & n28096;
  assign n28098 = ~n10074 & n28097;
  assign n28099 = ~n10780 & n28098;
  assign n28100 = n10640 & n28099;
  assign n28101 = n11323 & n28100;
  assign n28102 = n11342 & n28101;
  assign n28103 = ~n28095 & ~n28102;
  assign n28104 = n28085 & n28103;
  assign n28105 = n28054 & n28104;
  assign po109 = ~n27989 | ~n28105;
  assign n28107 = n4955 & n18694;
  assign n28108 = n7909 & n28107;
  assign n28109 = ~n2242 & n28108;
  assign n28110 = ~n3095 & n28109;
  assign n28111 = ~n3997 & n28110;
  assign n28112 = ~n4003 & n28111;
  assign n28113 = ~n4837 & n28112;
  assign n28114 = ~n5822 & n28113;
  assign n28115 = ~n6820 & n28114;
  assign n28116 = ~n7785 & n28115;
  assign n28117 = ~n9027 & n28116;
  assign n28118 = ~n10342 & n28117;
  assign n28119 = ~n10341 & n28118;
  assign n28120 = ~n10245 & n28119;
  assign n28121 = ~n10340 & n28120;
  assign n28122 = n10339 & n28121;
  assign n28123 = n10334 & n28122;
  assign n28124 = n10372 & n28123;
  assign n28125 = pi181 & ~n8900;
  assign n28126 = ~n10416 & n28125;
  assign n28127 = ~n9533 & n28126;
  assign n28128 = ~n10764 & n28127;
  assign n28129 = n10770 & n28128;
  assign n28130 = n10640 & n28129;
  assign n28131 = n10786 & n28130;
  assign n28132 = ~n28124 & ~n28131;
  assign n28133 = ~n8397 & n26211;
  assign n28134 = ~n10416 & n28133;
  assign n28135 = ~n10094 & n28134;
  assign n28136 = ~n10713 & n28135;
  assign n28137 = n10640 & n28136;
  assign n28138 = n11312 & n28137;
  assign n28139 = n11305 & n28138;
  assign n28140 = pi189 & ~n9687;
  assign n28141 = ~n9913 & n28140;
  assign n28142 = n11365 & n28141;
  assign n28143 = n9856 & n28142;
  assign n28144 = ~n9929 & n28143;
  assign n28145 = ~n10416 & n28144;
  assign n28146 = ~n10622 & n28145;
  assign n28147 = n10564 & n28146;
  assign n28148 = n11226 & n28147;
  assign n28149 = n11218 & n28148;
  assign n28150 = n11265 & n28149;
  assign n28151 = ~n28139 & ~n28150;
  assign n28152 = n28132 & n28151;
  assign n28153 = ~n9215 & n26113;
  assign n28154 = ~n10416 & n28153;
  assign n28155 = ~n10451 & n28154;
  assign n28156 = n10459 & n28155;
  assign n28157 = ~n9160 & n26084;
  assign n28158 = ~n10394 & n28157;
  assign n28159 = n10399 & n28158;
  assign n28160 = pi205 & ~n501;
  assign n28161 = n11440 & n28160;
  assign n28162 = n11446 & n28161;
  assign n28163 = n11437 & n28162;
  assign n28164 = ~n1172 & n28163;
  assign n28165 = ~n996 & n28164;
  assign n28166 = ~n2306 & n28165;
  assign n28167 = ~n500 & n28166;
  assign n28168 = n11004 & n28167;
  assign n28169 = n26550 & n28168;
  assign n28170 = n10980 & n28169;
  assign n28171 = n10971 & n28170;
  assign n28172 = n11172 & n28171;
  assign n28173 = ~n7236 & n28172;
  assign n28174 = ~n6137 & n28173;
  assign n28175 = n6193 & n28174;
  assign n28176 = n6134 & n28175;
  assign n28177 = ~n8867 & n28176;
  assign n28178 = ~n7235 & n28177;
  assign n28179 = n7296 & n28178;
  assign n28180 = n7231 & n28179;
  assign n28181 = ~n10027 & n28180;
  assign n28182 = ~n8866 & n28181;
  assign n28183 = n8898 & n28182;
  assign n28184 = n8863 & n28183;
  assign n28185 = ~n10026 & n28184;
  assign n28186 = n10072 & n28185;
  assign n28187 = n10021 & n28186;
  assign n28188 = pi213 & ~n501;
  assign n28189 = n26571 & n28188;
  assign n28190 = n26575 & n28189;
  assign n28191 = n11404 & n28190;
  assign n28192 = ~n1172 & n28191;
  assign n28193 = ~n996 & n28192;
  assign n28194 = ~n2306 & n28193;
  assign n28195 = ~n500 & n28194;
  assign n28196 = n10855 & n28195;
  assign n28197 = n26584 & n28196;
  assign n28198 = n10831 & n28197;
  assign n28199 = n10823 & n28198;
  assign n28200 = ~n7236 & n28199;
  assign n28201 = ~n6137 & n28200;
  assign n28202 = n6193 & n28201;
  assign n28203 = n6134 & n28202;
  assign n28204 = ~n8867 & n28203;
  assign n28205 = ~n7235 & n28204;
  assign n28206 = n7296 & n28205;
  assign n28207 = n7231 & n28206;
  assign n28208 = ~n10027 & n28207;
  assign n28209 = ~n8866 & n28208;
  assign n28210 = n8898 & n28209;
  assign n28211 = n8863 & n28210;
  assign n28212 = ~n10788 & n28211;
  assign n28213 = ~n10026 & n28212;
  assign n28214 = n10072 & n28213;
  assign n28215 = n10021 & n28214;
  assign n28216 = ~n28187 & ~n28215;
  assign n28217 = ~n28159 & n28216;
  assign n28218 = ~n28156 & n28217;
  assign n28219 = ~n9307 & n26079;
  assign n28220 = ~n10416 & n28219;
  assign n28221 = ~n10452 & n28220;
  assign n28222 = n10552 & n28221;
  assign n28223 = n10546 & n28222;
  assign n28224 = ~n9381 & n26117;
  assign n28225 = ~n10416 & n28224;
  assign n28226 = n10564 & n28225;
  assign n28227 = n10627 & n28226;
  assign n28228 = n10621 & n28227;
  assign n28229 = ~n28223 & ~n28228;
  assign n28230 = n28218 & n28229;
  assign n28231 = n8363 & n26042;
  assign n28232 = ~n7869 & n28231;
  assign n28233 = ~n8346 & n28232;
  assign n28234 = ~n10714 & n28233;
  assign n28235 = ~n10416 & n28234;
  assign n28236 = ~n9485 & n28235;
  assign n28237 = ~n10713 & n28236;
  assign n28238 = n10640 & n28237;
  assign n28239 = n10712 & n28238;
  assign n28240 = n10740 & n28239;
  assign n28241 = n10602 & n21531;
  assign n28242 = ~n5808 & n28241;
  assign n28243 = ~n6056 & n28242;
  assign n28244 = ~n7073 & n28243;
  assign n28245 = ~n8179 & n28244;
  assign n28246 = ~n10568 & n28245;
  assign n28247 = ~n10416 & n28246;
  assign n28248 = ~n9344 & n28247;
  assign n28249 = ~n10567 & n28248;
  assign n28250 = n10566 & n28249;
  assign n28251 = n10563 & n28250;
  assign n28252 = n10593 & n28251;
  assign n28253 = ~n28240 & ~n28252;
  assign n28254 = n28230 & n28253;
  assign n28255 = n28152 & n28254;
  assign n28256 = ~n8291 & n26167;
  assign n28257 = ~n10416 & n28256;
  assign n28258 = ~n9453 & n28257;
  assign n28259 = ~n10696 & n28258;
  assign n28260 = n10702 & n28259;
  assign n28261 = n10640 & n28260;
  assign n28262 = n10695 & n28261;
  assign n28263 = pi045 & ~n1208;
  assign n28264 = n4920 & n28263;
  assign n28265 = n4931 & n28264;
  assign n28266 = n4928 & n28265;
  assign n28267 = ~n1372 & n28266;
  assign n28268 = ~n2243 & n28267;
  assign n28269 = ~n3104 & n28268;
  assign n28270 = ~n3971 & n28269;
  assign n28271 = ~n4003 & n28270;
  assign n28272 = ~n4872 & n28271;
  assign n28273 = ~n5801 & n28272;
  assign n28274 = ~n6739 & n28273;
  assign n28275 = ~n7807 & n28274;
  assign n28276 = ~n8989 & n28275;
  assign n28277 = ~n10293 & n28276;
  assign n28278 = ~n10292 & n28277;
  assign n28279 = ~n10273 & n28278;
  assign n28280 = ~n10291 & n28279;
  assign n28281 = n10290 & n28280;
  assign n28282 = n10285 & n28281;
  assign n28283 = n10326 & n28282;
  assign n28284 = ~n28262 & ~n28283;
  assign n28285 = n10376 & n26136;
  assign n28286 = n9115 & n28285;
  assign n28287 = ~n3066 & n28286;
  assign n28288 = ~n3983 & n28287;
  assign n28289 = ~n4003 & n28288;
  assign n28290 = ~n4024 & n28289;
  assign n28291 = ~n4999 & n28290;
  assign n28292 = ~n5827 & n28291;
  assign n28293 = ~n6893 & n28292;
  assign n28294 = ~n7890 & n28293;
  assign n28295 = ~n10206 & n28294;
  assign n28296 = ~n10205 & n28295;
  assign n28297 = ~n9131 & n28296;
  assign n28298 = ~n10204 & n28297;
  assign n28299 = n10203 & n28298;
  assign n28300 = n10198 & n28299;
  assign n28301 = n10277 & n28300;
  assign n28302 = pi093 & ~n3710;
  assign n28303 = n4096 & n28302;
  assign n28304 = n4104 & n28303;
  assign n28305 = n8056 & n28304;
  assign n28306 = ~n3940 & n28305;
  assign n28307 = ~n4001 & n28306;
  assign n28308 = ~n5043 & n28307;
  assign n28309 = ~n5943 & n28308;
  assign n28310 = ~n6951 & n28309;
  assign n28311 = ~n8037 & n28310;
  assign n28312 = ~n10417 & n28311;
  assign n28313 = ~n10416 & n28312;
  assign n28314 = ~n9200 & n28313;
  assign n28315 = ~n10415 & n28314;
  assign n28316 = n10414 & n28315;
  assign n28317 = n10409 & n28316;
  assign n28318 = n10444 & n28317;
  assign n28319 = ~n28301 & ~n28318;
  assign n28320 = n28284 & n28319;
  assign n28321 = pi141 & ~n6313;
  assign n28322 = n7169 & n28321;
  assign n28323 = n7177 & n28322;
  assign n28324 = n8261 & n28323;
  assign n28325 = ~n6784 & n28324;
  assign n28326 = ~n7158 & n28325;
  assign n28327 = ~n8250 & n28326;
  assign n28328 = ~n10642 & n28327;
  assign n28329 = ~n10416 & n28328;
  assign n28330 = ~n9414 & n28329;
  assign n28331 = ~n10641 & n28330;
  assign n28332 = n10640 & n28331;
  assign n28333 = n10638 & n28332;
  assign n28334 = n10666 & n28333;
  assign n28335 = pi109 & ~n4707;
  assign n28336 = n5083 & n28335;
  assign n28337 = n8096 & n28336;
  assign n28338 = n9263 & n28337;
  assign n28339 = ~n4817 & n28338;
  assign n28340 = ~n4902 & n28339;
  assign n28341 = ~n6001 & n28340;
  assign n28342 = ~n7014 & n28341;
  assign n28343 = ~n8114 & n28342;
  assign n28344 = ~n10496 & n28343;
  assign n28345 = ~n10416 & n28344;
  assign n28346 = ~n9276 & n28345;
  assign n28347 = ~n10495 & n28346;
  assign n28348 = n10494 & n28347;
  assign n28349 = n10490 & n28348;
  assign n28350 = n10522 & n28349;
  assign n28351 = ~n28334 & ~n28350;
  assign n28352 = n11378 & n26067;
  assign n28353 = n9942 & n28352;
  assign n28354 = ~n8834 & n28353;
  assign n28355 = ~n11273 & n28354;
  assign n28356 = ~n10416 & n28355;
  assign n28357 = ~n10002 & n28356;
  assign n28358 = ~n10780 & n28357;
  assign n28359 = n10640 & n28358;
  assign n28360 = n11272 & n28359;
  assign n28361 = n11296 & n28360;
  assign n28362 = pi197 & ~n11324;
  assign n28363 = ~n10416 & n28362;
  assign n28364 = ~n10074 & n28363;
  assign n28365 = ~n10780 & n28364;
  assign n28366 = n10640 & n28365;
  assign n28367 = n11323 & n28366;
  assign n28368 = n11342 & n28367;
  assign n28369 = ~n28361 & ~n28368;
  assign n28370 = n28351 & n28369;
  assign n28371 = n28320 & n28370;
  assign po110 = ~n28255 | ~n28371;
  assign n28373 = n4955 & n18732;
  assign n28374 = n7909 & n28373;
  assign n28375 = ~n2242 & n28374;
  assign n28376 = ~n3095 & n28375;
  assign n28377 = ~n3997 & n28376;
  assign n28378 = ~n4003 & n28377;
  assign n28379 = ~n4837 & n28378;
  assign n28380 = ~n5822 & n28379;
  assign n28381 = ~n6820 & n28380;
  assign n28382 = ~n7785 & n28381;
  assign n28383 = ~n9027 & n28382;
  assign n28384 = ~n10342 & n28383;
  assign n28385 = ~n10341 & n28384;
  assign n28386 = ~n10245 & n28385;
  assign n28387 = ~n10340 & n28386;
  assign n28388 = n10339 & n28387;
  assign n28389 = n10334 & n28388;
  assign n28390 = n10372 & n28389;
  assign n28391 = pi182 & ~n8900;
  assign n28392 = ~n10416 & n28391;
  assign n28393 = ~n9533 & n28392;
  assign n28394 = ~n10764 & n28393;
  assign n28395 = n10770 & n28394;
  assign n28396 = n10640 & n28395;
  assign n28397 = n10786 & n28396;
  assign n28398 = ~n28390 & ~n28397;
  assign n28399 = ~n8397 & n26444;
  assign n28400 = ~n10416 & n28399;
  assign n28401 = ~n10094 & n28400;
  assign n28402 = ~n10713 & n28401;
  assign n28403 = n10640 & n28402;
  assign n28404 = n11312 & n28403;
  assign n28405 = n11305 & n28404;
  assign n28406 = pi190 & ~n9687;
  assign n28407 = ~n9913 & n28406;
  assign n28408 = n11365 & n28407;
  assign n28409 = n9856 & n28408;
  assign n28410 = ~n9929 & n28409;
  assign n28411 = ~n10416 & n28410;
  assign n28412 = ~n10622 & n28411;
  assign n28413 = n10564 & n28412;
  assign n28414 = n11226 & n28413;
  assign n28415 = n11218 & n28414;
  assign n28416 = n11265 & n28415;
  assign n28417 = ~n28405 & ~n28416;
  assign n28418 = n28398 & n28417;
  assign n28419 = ~n9215 & n26346;
  assign n28420 = ~n10416 & n28419;
  assign n28421 = ~n10451 & n28420;
  assign n28422 = n10459 & n28421;
  assign n28423 = ~n9160 & n26317;
  assign n28424 = ~n10394 & n28423;
  assign n28425 = n10399 & n28424;
  assign n28426 = pi206 & ~n501;
  assign n28427 = n11440 & n28426;
  assign n28428 = n11446 & n28427;
  assign n28429 = n11437 & n28428;
  assign n28430 = ~n1172 & n28429;
  assign n28431 = ~n996 & n28430;
  assign n28432 = ~n2306 & n28431;
  assign n28433 = ~n500 & n28432;
  assign n28434 = n11004 & n28433;
  assign n28435 = n26550 & n28434;
  assign n28436 = n10980 & n28435;
  assign n28437 = n10971 & n28436;
  assign n28438 = n11172 & n28437;
  assign n28439 = ~n7236 & n28438;
  assign n28440 = ~n6137 & n28439;
  assign n28441 = n6193 & n28440;
  assign n28442 = n6134 & n28441;
  assign n28443 = ~n8867 & n28442;
  assign n28444 = ~n7235 & n28443;
  assign n28445 = n7296 & n28444;
  assign n28446 = n7231 & n28445;
  assign n28447 = ~n10027 & n28446;
  assign n28448 = ~n8866 & n28447;
  assign n28449 = n8898 & n28448;
  assign n28450 = n8863 & n28449;
  assign n28451 = ~n10026 & n28450;
  assign n28452 = n10072 & n28451;
  assign n28453 = n10021 & n28452;
  assign n28454 = pi214 & ~n501;
  assign n28455 = n26571 & n28454;
  assign n28456 = n26575 & n28455;
  assign n28457 = n11404 & n28456;
  assign n28458 = ~n1172 & n28457;
  assign n28459 = ~n996 & n28458;
  assign n28460 = ~n2306 & n28459;
  assign n28461 = ~n500 & n28460;
  assign n28462 = n10855 & n28461;
  assign n28463 = n26584 & n28462;
  assign n28464 = n10831 & n28463;
  assign n28465 = n10823 & n28464;
  assign n28466 = ~n7236 & n28465;
  assign n28467 = ~n6137 & n28466;
  assign n28468 = n6193 & n28467;
  assign n28469 = n6134 & n28468;
  assign n28470 = ~n8867 & n28469;
  assign n28471 = ~n7235 & n28470;
  assign n28472 = n7296 & n28471;
  assign n28473 = n7231 & n28472;
  assign n28474 = ~n10027 & n28473;
  assign n28475 = ~n8866 & n28474;
  assign n28476 = n8898 & n28475;
  assign n28477 = n8863 & n28476;
  assign n28478 = ~n10788 & n28477;
  assign n28479 = ~n10026 & n28478;
  assign n28480 = n10072 & n28479;
  assign n28481 = n10021 & n28480;
  assign n28482 = ~n28453 & ~n28481;
  assign n28483 = ~n28425 & n28482;
  assign n28484 = ~n28422 & n28483;
  assign n28485 = ~n9307 & n26312;
  assign n28486 = ~n10416 & n28485;
  assign n28487 = ~n10452 & n28486;
  assign n28488 = n10552 & n28487;
  assign n28489 = n10546 & n28488;
  assign n28490 = ~n9381 & n26350;
  assign n28491 = ~n10416 & n28490;
  assign n28492 = n10564 & n28491;
  assign n28493 = n10627 & n28492;
  assign n28494 = n10621 & n28493;
  assign n28495 = ~n28489 & ~n28494;
  assign n28496 = n28484 & n28495;
  assign n28497 = n8363 & n26275;
  assign n28498 = ~n7869 & n28497;
  assign n28499 = ~n8346 & n28498;
  assign n28500 = ~n10714 & n28499;
  assign n28501 = ~n10416 & n28500;
  assign n28502 = ~n9485 & n28501;
  assign n28503 = ~n10713 & n28502;
  assign n28504 = n10640 & n28503;
  assign n28505 = n10712 & n28504;
  assign n28506 = n10740 & n28505;
  assign n28507 = n10602 & n21657;
  assign n28508 = ~n5808 & n28507;
  assign n28509 = ~n6056 & n28508;
  assign n28510 = ~n7073 & n28509;
  assign n28511 = ~n8179 & n28510;
  assign n28512 = ~n10568 & n28511;
  assign n28513 = ~n10416 & n28512;
  assign n28514 = ~n9344 & n28513;
  assign n28515 = ~n10567 & n28514;
  assign n28516 = n10566 & n28515;
  assign n28517 = n10563 & n28516;
  assign n28518 = n10593 & n28517;
  assign n28519 = ~n28506 & ~n28518;
  assign n28520 = n28496 & n28519;
  assign n28521 = n28418 & n28520;
  assign n28522 = ~n8291 & n26400;
  assign n28523 = ~n10416 & n28522;
  assign n28524 = ~n9453 & n28523;
  assign n28525 = ~n10696 & n28524;
  assign n28526 = n10702 & n28525;
  assign n28527 = n10640 & n28526;
  assign n28528 = n10695 & n28527;
  assign n28529 = pi046 & ~n1208;
  assign n28530 = n4920 & n28529;
  assign n28531 = n4931 & n28530;
  assign n28532 = n4928 & n28531;
  assign n28533 = ~n1372 & n28532;
  assign n28534 = ~n2243 & n28533;
  assign n28535 = ~n3104 & n28534;
  assign n28536 = ~n3971 & n28535;
  assign n28537 = ~n4003 & n28536;
  assign n28538 = ~n4872 & n28537;
  assign n28539 = ~n5801 & n28538;
  assign n28540 = ~n6739 & n28539;
  assign n28541 = ~n7807 & n28540;
  assign n28542 = ~n8989 & n28541;
  assign n28543 = ~n10293 & n28542;
  assign n28544 = ~n10292 & n28543;
  assign n28545 = ~n10273 & n28544;
  assign n28546 = ~n10291 & n28545;
  assign n28547 = n10290 & n28546;
  assign n28548 = n10285 & n28547;
  assign n28549 = n10326 & n28548;
  assign n28550 = ~n28528 & ~n28549;
  assign n28551 = n10376 & n26369;
  assign n28552 = n9115 & n28551;
  assign n28553 = ~n3066 & n28552;
  assign n28554 = ~n3983 & n28553;
  assign n28555 = ~n4003 & n28554;
  assign n28556 = ~n4024 & n28555;
  assign n28557 = ~n4999 & n28556;
  assign n28558 = ~n5827 & n28557;
  assign n28559 = ~n6893 & n28558;
  assign n28560 = ~n7890 & n28559;
  assign n28561 = ~n10206 & n28560;
  assign n28562 = ~n10205 & n28561;
  assign n28563 = ~n9131 & n28562;
  assign n28564 = ~n10204 & n28563;
  assign n28565 = n10203 & n28564;
  assign n28566 = n10198 & n28565;
  assign n28567 = n10277 & n28566;
  assign n28568 = pi094 & ~n3710;
  assign n28569 = n4096 & n28568;
  assign n28570 = n4104 & n28569;
  assign n28571 = n8056 & n28570;
  assign n28572 = ~n3940 & n28571;
  assign n28573 = ~n4001 & n28572;
  assign n28574 = ~n5043 & n28573;
  assign n28575 = ~n5943 & n28574;
  assign n28576 = ~n6951 & n28575;
  assign n28577 = ~n8037 & n28576;
  assign n28578 = ~n10417 & n28577;
  assign n28579 = ~n10416 & n28578;
  assign n28580 = ~n9200 & n28579;
  assign n28581 = ~n10415 & n28580;
  assign n28582 = n10414 & n28581;
  assign n28583 = n10409 & n28582;
  assign n28584 = n10444 & n28583;
  assign n28585 = ~n28567 & ~n28584;
  assign n28586 = n28550 & n28585;
  assign n28587 = pi142 & ~n6313;
  assign n28588 = n7169 & n28587;
  assign n28589 = n7177 & n28588;
  assign n28590 = n8261 & n28589;
  assign n28591 = ~n6784 & n28590;
  assign n28592 = ~n7158 & n28591;
  assign n28593 = ~n8250 & n28592;
  assign n28594 = ~n10642 & n28593;
  assign n28595 = ~n10416 & n28594;
  assign n28596 = ~n9414 & n28595;
  assign n28597 = ~n10641 & n28596;
  assign n28598 = n10640 & n28597;
  assign n28599 = n10638 & n28598;
  assign n28600 = n10666 & n28599;
  assign n28601 = pi110 & ~n4707;
  assign n28602 = n5083 & n28601;
  assign n28603 = n8096 & n28602;
  assign n28604 = n9263 & n28603;
  assign n28605 = ~n4817 & n28604;
  assign n28606 = ~n4902 & n28605;
  assign n28607 = ~n6001 & n28606;
  assign n28608 = ~n7014 & n28607;
  assign n28609 = ~n8114 & n28608;
  assign n28610 = ~n10496 & n28609;
  assign n28611 = ~n10416 & n28610;
  assign n28612 = ~n9276 & n28611;
  assign n28613 = ~n10495 & n28612;
  assign n28614 = n10494 & n28613;
  assign n28615 = n10490 & n28614;
  assign n28616 = n10522 & n28615;
  assign n28617 = ~n28600 & ~n28616;
  assign n28618 = n11378 & n26300;
  assign n28619 = n9942 & n28618;
  assign n28620 = ~n8834 & n28619;
  assign n28621 = ~n11273 & n28620;
  assign n28622 = ~n10416 & n28621;
  assign n28623 = ~n10002 & n28622;
  assign n28624 = ~n10780 & n28623;
  assign n28625 = n10640 & n28624;
  assign n28626 = n11272 & n28625;
  assign n28627 = n11296 & n28626;
  assign n28628 = pi198 & ~n11324;
  assign n28629 = ~n10416 & n28628;
  assign n28630 = ~n10074 & n28629;
  assign n28631 = ~n10780 & n28630;
  assign n28632 = n10640 & n28631;
  assign n28633 = n11323 & n28632;
  assign n28634 = n11342 & n28633;
  assign n28635 = ~n28627 & ~n28634;
  assign n28636 = n28617 & n28635;
  assign n28637 = n28586 & n28636;
  assign po111 = ~n28521 | ~n28637;
  assign n28639 = ~n10554 & n26612;
  assign n28640 = ~n11510 & n28639;
  assign n28641 = ~n11506 & n28640;
  assign n28642 = n11957 & n28641;
  assign n28643 = n11952 & n28642;
  assign n28644 = ~n10400 & n26536;
  assign n28645 = ~n11790 & n28644;
  assign n28646 = n11795 & n28645;
  assign n28647 = ~n1493 & ~n9651;
  assign n28648 = n12496 & n28647;
  assign n28649 = n14227 & n28648;
  assign n28650 = n12535 & n28649;
  assign n28651 = n12549 & n14210;
  assign n28652 = n12604 & n28651;
  assign n28653 = n11402 & n18073;
  assign n28654 = n28652 & n28653;
  assign n28655 = pi223 & ~n501;
  assign n28656 = n12872 & n28655;
  assign n28657 = n14253 & n28656;
  assign n28658 = n12564 & n28657;
  assign n28659 = n28654 & n28658;
  assign n28660 = n12548 & n28659;
  assign n28661 = ~n1172 & n28660;
  assign n28662 = ~n996 & n28661;
  assign n28663 = ~n2306 & n28662;
  assign n28664 = n12571 & n28663;
  assign n28665 = n6677 & n28664;
  assign n28666 = n12580 & n28665;
  assign n28667 = n3822 & n12498;
  assign n28668 = n12583 & n28667;
  assign n28669 = n28666 & n28668;
  assign n28670 = n12542 & n28669;
  assign n28671 = n28650 & n28670;
  assign n28672 = ~n7236 & n28671;
  assign n28673 = ~n6137 & n28672;
  assign n28674 = n6193 & n28673;
  assign n28675 = n6134 & n28674;
  assign n28676 = ~n8867 & n28675;
  assign n28677 = ~n7235 & n28676;
  assign n28678 = n7296 & n28677;
  assign n28679 = n7231 & n28678;
  assign n28680 = ~n10027 & n28679;
  assign n28681 = ~n8866 & n28680;
  assign n28682 = n8898 & n28681;
  assign n28683 = n8863 & n28682;
  assign n28684 = ~n2726 & ~n3770;
  assign n28685 = n14210 & n28684;
  assign n28686 = n12604 & n28685;
  assign n28687 = n12607 & n15998;
  assign n28688 = n11402 & n28687;
  assign n28689 = n28686 & n28688;
  assign n28690 = pi215 & ~n501;
  assign n28691 = n12611 & n28690;
  assign n28692 = n26571 & n28691;
  assign n28693 = n12619 & n28692;
  assign n28694 = n28689 & n28693;
  assign n28695 = n12601 & n28694;
  assign n28696 = ~n1172 & n28695;
  assign n28697 = ~n996 & n28696;
  assign n28698 = ~n2306 & n28697;
  assign n28699 = n12626 & n28698;
  assign n28700 = n12628 & n28699;
  assign n28701 = n3823 & n28700;
  assign n28702 = n12634 & n28701;
  assign n28703 = n12682 & n28702;
  assign n28704 = n12844 & n28703;
  assign n28705 = ~n7236 & n28704;
  assign n28706 = ~n6137 & n28705;
  assign n28707 = n6193 & n28706;
  assign n28708 = n6134 & n28707;
  assign n28709 = ~n8867 & n28708;
  assign n28710 = ~n7235 & n28709;
  assign n28711 = n7296 & n28710;
  assign n28712 = n7231 & n28711;
  assign n28713 = ~n10027 & n28712;
  assign n28714 = ~n8866 & n28713;
  assign n28715 = n8898 & n28714;
  assign n28716 = n8863 & n28715;
  assign n28717 = ~n28683 & ~n28716;
  assign n28718 = ~n10788 & ~n28717;
  assign n28719 = ~n10026 & n28718;
  assign n28720 = n10072 & n28719;
  assign n28721 = n10021 & n28720;
  assign n28722 = ~n28646 & ~n28721;
  assign n28723 = ~n28643 & n28722;
  assign n28724 = ~n10629 & n26607;
  assign n28725 = ~n11510 & n28724;
  assign n28726 = n11970 & n28725;
  assign n28727 = n12039 & n28726;
  assign n28728 = n12034 & n28727;
  assign n28729 = ~n10460 & n26532;
  assign n28730 = ~n11510 & n28729;
  assign n28731 = ~n11852 & n28730;
  assign n28732 = n11859 & n28731;
  assign n28733 = ~n28728 & ~n28732;
  assign n28734 = n28723 & n28733;
  assign n28735 = ~n8574 & n24608;
  assign n28736 = n9934 & n28735;
  assign n28737 = n8545 & n28736;
  assign n28738 = ~n8834 & n28737;
  assign n28739 = ~n10002 & n28738;
  assign n28740 = ~n12212 & n28739;
  assign n28741 = ~n12211 & n28740;
  assign n28742 = ~n11510 & n28741;
  assign n28743 = ~n11297 & n28742;
  assign n28744 = ~n11478 & n28743;
  assign n28745 = n11508 & n28744;
  assign n28746 = n12210 & n28745;
  assign n28747 = n12239 & n28746;
  assign n28748 = n2784 & n3852;
  assign n28749 = n23168 & n28748;
  assign n28750 = ~n3066 & n28749;
  assign n28751 = ~n3983 & n28750;
  assign n28752 = ~n4003 & n28751;
  assign n28753 = ~n4024 & n28752;
  assign n28754 = ~n4999 & n28753;
  assign n28755 = ~n5827 & n28754;
  assign n28756 = ~n6893 & n28755;
  assign n28757 = ~n7890 & n28756;
  assign n28758 = ~n9131 & n28757;
  assign n28759 = ~n11627 & n28758;
  assign n28760 = ~n11626 & n28759;
  assign n28761 = ~n11625 & n28760;
  assign n28762 = ~n10278 & n28761;
  assign n28763 = ~n11624 & n28762;
  assign n28764 = n11623 & n28763;
  assign n28765 = n11618 & n28764;
  assign n28766 = n11661 & n28765;
  assign n28767 = ~n28747 & ~n28766;
  assign n28768 = pi191 & ~n10074;
  assign n28769 = ~n11510 & n28768;
  assign n28770 = ~n11343 & n28769;
  assign n28771 = ~n11509 & n28770;
  assign n28772 = n11508 & n28771;
  assign n28773 = n11503 & n28772;
  assign n28774 = n11550 & n28773;
  assign n28775 = n7175 & n26737;
  assign n28776 = n26733 & n28775;
  assign n28777 = ~n6784 & n28776;
  assign n28778 = ~n7158 & n28777;
  assign n28779 = ~n8250 & n28778;
  assign n28780 = ~n9414 & n28779;
  assign n28781 = ~n12053 & n28780;
  assign n28782 = ~n12052 & n28781;
  assign n28783 = ~n11510 & n28782;
  assign n28784 = ~n10667 & n28783;
  assign n28785 = ~n12051 & n28784;
  assign n28786 = n11508 & n28785;
  assign n28787 = n12050 & n28786;
  assign n28788 = n12082 & n28787;
  assign n28789 = ~n28774 & ~n28788;
  assign n28790 = n28767 & n28789;
  assign n28791 = n28734 & n28790;
  assign n28792 = ~n9453 & n26658;
  assign n28793 = ~n11510 & n28792;
  assign n28794 = ~n10705 & n28793;
  assign n28795 = ~n12112 & n28794;
  assign n28796 = n12118 & n28795;
  assign n28797 = n11508 & n28796;
  assign n28798 = n12111 & n28797;
  assign n28799 = pi207 & ~n10879;
  assign n28800 = ~n12412 & n28799;
  assign n28801 = ~n11510 & n28800;
  assign n28802 = ~n11505 & n28801;
  assign n28803 = n11970 & n28802;
  assign n28804 = n12325 & n28803;
  assign n28805 = n12411 & n28804;
  assign n28806 = n12470 & n28805;
  assign n28807 = ~n28798 & ~n28806;
  assign n28808 = ~n9533 & n26651;
  assign n28809 = ~n11510 & n28808;
  assign n28810 = ~n10787 & n28809;
  assign n28811 = ~n11478 & n28810;
  assign n28812 = n11593 & n28811;
  assign n28813 = n11508 & n28812;
  assign n28814 = n11610 & n28813;
  assign n28815 = pi055 & ~n2172;
  assign n28816 = ~n2173 & n28815;
  assign n28817 = ~n2171 & n28816;
  assign n28818 = ~n1679 & n28817;
  assign n28819 = n1741 & n28818;
  assign n28820 = n1619 & n28819;
  assign n28821 = ~n2242 & n28820;
  assign n28822 = ~n3095 & n28821;
  assign n28823 = ~n3997 & n28822;
  assign n28824 = ~n4003 & n28823;
  assign n28825 = ~n4837 & n28824;
  assign n28826 = ~n5822 & n28825;
  assign n28827 = ~n6820 & n28826;
  assign n28828 = ~n7785 & n28827;
  assign n28829 = ~n9027 & n28828;
  assign n28830 = ~n10245 & n28829;
  assign n28831 = ~n11733 & n28830;
  assign n28832 = ~n11732 & n28831;
  assign n28833 = ~n11731 & n28832;
  assign n28834 = ~n11536 & n28833;
  assign n28835 = ~n11730 & n28834;
  assign n28836 = n11729 & n28835;
  assign n28837 = n11724 & n28836;
  assign n28838 = n11768 & n28837;
  assign n28839 = ~n28814 & ~n28838;
  assign n28840 = n28807 & n28839;
  assign n28841 = ~n10094 & n26666;
  assign n28842 = ~n11510 & n28841;
  assign n28843 = ~n11318 & n28842;
  assign n28844 = ~n11501 & n28843;
  assign n28845 = n11508 & n28844;
  assign n28846 = n12175 & n28845;
  assign n28847 = n12168 & n28846;
  assign n28848 = pi183 & ~n9687;
  assign n28849 = n12275 & n28848;
  assign n28850 = n11562 & n28849;
  assign n28851 = n11560 & n28850;
  assign n28852 = ~n9929 & n28851;
  assign n28853 = ~n11558 & n28852;
  assign n28854 = ~n11557 & n28853;
  assign n28855 = ~n11510 & n28854;
  assign n28856 = ~n11266 & n28855;
  assign n28857 = ~n11509 & n28856;
  assign n28858 = n11508 & n28857;
  assign n28859 = n11556 & n28858;
  assign n28860 = n11587 & n28859;
  assign n28861 = ~n28847 & ~n28860;
  assign n28862 = pi087 & ~n3399;
  assign n28863 = ~n3400 & n28862;
  assign n28864 = ~n3398 & n28863;
  assign n28865 = ~n3710 & n28864;
  assign n28866 = n4096 & n28865;
  assign n28867 = n4104 & n28866;
  assign n28868 = ~n3940 & n28867;
  assign n28869 = ~n4001 & n28868;
  assign n28870 = ~n5043 & n28869;
  assign n28871 = ~n5943 & n28870;
  assign n28872 = ~n6951 & n28871;
  assign n28873 = ~n8037 & n28872;
  assign n28874 = ~n9200 & n28873;
  assign n28875 = ~n11813 & n28874;
  assign n28876 = ~n11812 & n28875;
  assign n28877 = ~n11510 & n28876;
  assign n28878 = ~n10445 & n28877;
  assign n28879 = ~n11811 & n28878;
  assign n28880 = n11810 & n28879;
  assign n28881 = n11805 & n28880;
  assign n28882 = n11845 & n28881;
  assign n28883 = n5084 & n26510;
  assign n28884 = n5083 & n26515;
  assign n28885 = n28883 & n28884;
  assign n28886 = ~n4817 & n28885;
  assign n28887 = ~n4902 & n28886;
  assign n28888 = ~n6001 & n28887;
  assign n28889 = ~n7014 & n28888;
  assign n28890 = ~n8114 & n28889;
  assign n28891 = ~n9276 & n28890;
  assign n28892 = ~n11898 & n28891;
  assign n28893 = ~n11897 & n28892;
  assign n28894 = ~n11510 & n28893;
  assign n28895 = ~n10523 & n28894;
  assign n28896 = ~n11896 & n28895;
  assign n28897 = n11895 & n28896;
  assign n28898 = n11891 & n28897;
  assign n28899 = n11927 & n28898;
  assign n28900 = ~n28882 & ~n28899;
  assign n28901 = n28861 & n28900;
  assign n28902 = ~n718 & ~n841;
  assign n28903 = n13201 & n28902;
  assign n28904 = pi039 & ~n807;
  assign n28905 = ~n808 & n28904;
  assign n28906 = ~n806 & n28905;
  assign n28907 = ~n1208 & n28906;
  assign n28908 = n4920 & n28907;
  assign n28909 = n28903 & n28908;
  assign n28910 = ~n1372 & n28909;
  assign n28911 = ~n2243 & n28910;
  assign n28912 = ~n3104 & n28911;
  assign n28913 = ~n3971 & n28912;
  assign n28914 = ~n4003 & n28913;
  assign n28915 = ~n4872 & n28914;
  assign n28916 = ~n5801 & n28915;
  assign n28917 = ~n6739 & n28916;
  assign n28918 = ~n7807 & n28917;
  assign n28919 = ~n8989 & n28918;
  assign n28920 = ~n10273 & n28919;
  assign n28921 = ~n11678 & n28920;
  assign n28922 = ~n11677 & n28921;
  assign n28923 = ~n11676 & n28922;
  assign n28924 = ~n11499 & n28923;
  assign n28925 = ~n11675 & n28924;
  assign n28926 = n11674 & n28925;
  assign n28927 = n11669 & n28926;
  assign n28928 = n11716 & n28927;
  assign n28929 = n7096 & n26619;
  assign n28930 = n12013 & n28929;
  assign n28931 = ~n5808 & n28930;
  assign n28932 = ~n6056 & n28931;
  assign n28933 = ~n7073 & n28932;
  assign n28934 = ~n8179 & n28933;
  assign n28935 = ~n9344 & n28934;
  assign n28936 = ~n11974 & n28935;
  assign n28937 = ~n11973 & n28936;
  assign n28938 = ~n11510 & n28937;
  assign n28939 = ~n10594 & n28938;
  assign n28940 = ~n11972 & n28939;
  assign n28941 = n11971 & n28940;
  assign n28942 = n11968 & n28941;
  assign n28943 = n12004 & n28942;
  assign n28944 = ~n28928 & ~n28943;
  assign n28945 = n12131 & n23137;
  assign n28946 = ~n7869 & n28945;
  assign n28947 = ~n8346 & n28946;
  assign n28948 = ~n9485 & n28947;
  assign n28949 = ~n12130 & n28948;
  assign n28950 = ~n12129 & n28949;
  assign n28951 = ~n11510 & n28950;
  assign n28952 = ~n10741 & n28951;
  assign n28953 = ~n11501 & n28952;
  assign n28954 = n11508 & n28953;
  assign n28955 = n12128 & n28954;
  assign n28956 = n12157 & n28955;
  assign n28957 = pi199 & ~n10939;
  assign n28958 = n12473 & n28957;
  assign n28959 = n12317 & n28958;
  assign n28960 = n12316 & n28959;
  assign n28961 = ~n11188 & n28960;
  assign n28962 = ~n12314 & n28961;
  assign n28963 = ~n11510 & n28962;
  assign n28964 = ~n11505 & n28963;
  assign n28965 = n11970 & n28964;
  assign n28966 = n12325 & n28965;
  assign n28967 = n12313 & n28966;
  assign n28968 = n12379 & n28967;
  assign n28969 = ~n28956 & ~n28968;
  assign n28970 = n28944 & n28969;
  assign n28971 = n28901 & n28970;
  assign n28972 = n28840 & n28971;
  assign po112 = ~n28791 | ~n28972;
  assign n28974 = ~n10460 & n26833;
  assign n28975 = ~n11510 & n28974;
  assign n28976 = ~n11852 & n28975;
  assign n28977 = n11859 & n28976;
  assign n28978 = ~n10400 & n26837;
  assign n28979 = ~n11790 & n28978;
  assign n28980 = n11795 & n28979;
  assign n28981 = pi224 & ~n501;
  assign n28982 = n12872 & n28981;
  assign n28983 = n14253 & n28982;
  assign n28984 = n12564 & n28983;
  assign n28985 = n28654 & n28984;
  assign n28986 = n12548 & n28985;
  assign n28987 = ~n1172 & n28986;
  assign n28988 = ~n996 & n28987;
  assign n28989 = ~n2306 & n28988;
  assign n28990 = n12571 & n28989;
  assign n28991 = n6677 & n28990;
  assign n28992 = n12580 & n28991;
  assign n28993 = n28668 & n28992;
  assign n28994 = n12542 & n28993;
  assign n28995 = n28650 & n28994;
  assign n28996 = ~n7236 & n28995;
  assign n28997 = ~n6137 & n28996;
  assign n28998 = n6193 & n28997;
  assign n28999 = n6134 & n28998;
  assign n29000 = ~n8867 & n28999;
  assign n29001 = ~n7235 & n29000;
  assign n29002 = n7296 & n29001;
  assign n29003 = n7231 & n29002;
  assign n29004 = ~n10027 & n29003;
  assign n29005 = ~n8866 & n29004;
  assign n29006 = n8898 & n29005;
  assign n29007 = n8863 & n29006;
  assign n29008 = pi216 & ~n501;
  assign n29009 = n12611 & n29008;
  assign n29010 = n26571 & n29009;
  assign n29011 = n12619 & n29010;
  assign n29012 = n28689 & n29011;
  assign n29013 = n12601 & n29012;
  assign n29014 = ~n1172 & n29013;
  assign n29015 = ~n996 & n29014;
  assign n29016 = ~n2306 & n29015;
  assign n29017 = n12626 & n29016;
  assign n29018 = n12628 & n29017;
  assign n29019 = n3823 & n29018;
  assign n29020 = n12634 & n29019;
  assign n29021 = n12682 & n29020;
  assign n29022 = n12844 & n29021;
  assign n29023 = ~n7236 & n29022;
  assign n29024 = ~n6137 & n29023;
  assign n29025 = n6193 & n29024;
  assign n29026 = n6134 & n29025;
  assign n29027 = ~n8867 & n29026;
  assign n29028 = ~n7235 & n29027;
  assign n29029 = n7296 & n29028;
  assign n29030 = n7231 & n29029;
  assign n29031 = ~n10027 & n29030;
  assign n29032 = ~n8866 & n29031;
  assign n29033 = n8898 & n29032;
  assign n29034 = n8863 & n29033;
  assign n29035 = ~n29007 & ~n29034;
  assign n29036 = ~n10788 & ~n29035;
  assign n29037 = ~n10026 & n29036;
  assign n29038 = n10072 & n29037;
  assign n29039 = n10021 & n29038;
  assign n29040 = ~n28980 & ~n29039;
  assign n29041 = ~n28977 & n29040;
  assign n29042 = ~n10554 & n26899;
  assign n29043 = ~n11510 & n29042;
  assign n29044 = ~n11506 & n29043;
  assign n29045 = n11957 & n29044;
  assign n29046 = n11952 & n29045;
  assign n29047 = ~n10629 & n26904;
  assign n29048 = ~n11510 & n29047;
  assign n29049 = n11970 & n29048;
  assign n29050 = n12039 & n29049;
  assign n29051 = n12034 & n29050;
  assign n29052 = ~n29046 & ~n29051;
  assign n29053 = n29041 & n29052;
  assign n29054 = n7177 & n27007;
  assign n29055 = n8261 & n29054;
  assign n29056 = ~n6784 & n29055;
  assign n29057 = ~n7158 & n29056;
  assign n29058 = ~n8250 & n29057;
  assign n29059 = ~n9414 & n29058;
  assign n29060 = ~n12053 & n29059;
  assign n29061 = ~n12052 & n29060;
  assign n29062 = ~n11510 & n29061;
  assign n29063 = ~n10667 & n29062;
  assign n29064 = ~n12051 & n29063;
  assign n29065 = n11508 & n29064;
  assign n29066 = n12050 & n29065;
  assign n29067 = n12082 & n29066;
  assign n29068 = n11681 & n26952;
  assign n29069 = n11680 & n29068;
  assign n29070 = ~n1372 & n29069;
  assign n29071 = ~n2243 & n29070;
  assign n29072 = ~n3104 & n29071;
  assign n29073 = ~n3971 & n29072;
  assign n29074 = ~n4003 & n29073;
  assign n29075 = ~n4872 & n29074;
  assign n29076 = ~n5801 & n29075;
  assign n29077 = ~n6739 & n29076;
  assign n29078 = ~n7807 & n29077;
  assign n29079 = ~n8989 & n29078;
  assign n29080 = ~n10273 & n29079;
  assign n29081 = ~n11678 & n29080;
  assign n29082 = ~n11677 & n29081;
  assign n29083 = ~n11676 & n29082;
  assign n29084 = ~n11499 & n29083;
  assign n29085 = ~n11675 & n29084;
  assign n29086 = n11674 & n29085;
  assign n29087 = n11669 & n29086;
  assign n29088 = n11716 & n29087;
  assign n29089 = ~n29067 & ~n29088;
  assign n29090 = n5062 & n26787;
  assign n29091 = n11861 & n29090;
  assign n29092 = ~n3940 & n29091;
  assign n29093 = ~n4001 & n29092;
  assign n29094 = ~n5043 & n29093;
  assign n29095 = ~n5943 & n29094;
  assign n29096 = ~n6951 & n29095;
  assign n29097 = ~n8037 & n29096;
  assign n29098 = ~n9200 & n29097;
  assign n29099 = ~n11813 & n29098;
  assign n29100 = ~n11812 & n29099;
  assign n29101 = ~n11510 & n29100;
  assign n29102 = ~n10445 & n29101;
  assign n29103 = ~n11811 & n29102;
  assign n29104 = n11810 & n29103;
  assign n29105 = n11805 & n29104;
  assign n29106 = n11845 & n29105;
  assign n29107 = ~n9533 & n26944;
  assign n29108 = ~n11510 & n29107;
  assign n29109 = ~n10787 & n29108;
  assign n29110 = ~n11478 & n29109;
  assign n29111 = n11593 & n29110;
  assign n29112 = n11508 & n29111;
  assign n29113 = n11610 & n29112;
  assign n29114 = ~n29106 & ~n29113;
  assign n29115 = n29089 & n29114;
  assign n29116 = n29053 & n29115;
  assign n29117 = n12182 & n23404;
  assign n29118 = ~n7869 & n29117;
  assign n29119 = ~n8346 & n29118;
  assign n29120 = ~n9485 & n29119;
  assign n29121 = ~n12130 & n29120;
  assign n29122 = ~n12129 & n29121;
  assign n29123 = ~n11510 & n29122;
  assign n29124 = ~n10741 & n29123;
  assign n29125 = ~n11501 & n29124;
  assign n29126 = n11508 & n29125;
  assign n29127 = n12128 & n29126;
  assign n29128 = n12157 & n29127;
  assign n29129 = ~n10094 & n26973;
  assign n29130 = ~n11510 & n29129;
  assign n29131 = ~n11318 & n29130;
  assign n29132 = ~n11501 & n29131;
  assign n29133 = n11508 & n29132;
  assign n29134 = n12175 & n29133;
  assign n29135 = n12168 & n29134;
  assign n29136 = ~n29128 & ~n29135;
  assign n29137 = n11378 & n24970;
  assign n29138 = n9942 & n29137;
  assign n29139 = ~n8834 & n29138;
  assign n29140 = ~n10002 & n29139;
  assign n29141 = ~n12212 & n29140;
  assign n29142 = ~n12211 & n29141;
  assign n29143 = ~n11510 & n29142;
  assign n29144 = ~n11297 & n29143;
  assign n29145 = ~n11478 & n29144;
  assign n29146 = n11508 & n29145;
  assign n29147 = n12210 & n29146;
  assign n29148 = n12239 & n29147;
  assign n29149 = n9115 & n21884;
  assign n29150 = ~n3066 & n29149;
  assign n29151 = ~n3983 & n29150;
  assign n29152 = ~n4003 & n29151;
  assign n29153 = ~n4024 & n29152;
  assign n29154 = ~n4999 & n29153;
  assign n29155 = ~n5827 & n29154;
  assign n29156 = ~n6893 & n29155;
  assign n29157 = ~n7890 & n29156;
  assign n29158 = ~n9131 & n29157;
  assign n29159 = ~n11627 & n29158;
  assign n29160 = ~n11626 & n29159;
  assign n29161 = ~n11625 & n29160;
  assign n29162 = ~n10278 & n29161;
  assign n29163 = ~n11624 & n29162;
  assign n29164 = n11623 & n29163;
  assign n29165 = n11618 & n29164;
  assign n29166 = n11661 & n29165;
  assign n29167 = ~n29148 & ~n29166;
  assign n29168 = n29136 & n29167;
  assign n29169 = pi208 & ~n10879;
  assign n29170 = ~n12412 & n29169;
  assign n29171 = ~n11510 & n29170;
  assign n29172 = ~n11505 & n29171;
  assign n29173 = n11970 & n29172;
  assign n29174 = n12325 & n29173;
  assign n29175 = n12411 & n29174;
  assign n29176 = n12470 & n29175;
  assign n29177 = n5085 & n26815;
  assign n29178 = n11931 & n29177;
  assign n29179 = ~n4817 & n29178;
  assign n29180 = ~n4902 & n29179;
  assign n29181 = ~n6001 & n29180;
  assign n29182 = ~n7014 & n29181;
  assign n29183 = ~n8114 & n29182;
  assign n29184 = ~n9276 & n29183;
  assign n29185 = ~n11898 & n29184;
  assign n29186 = ~n11897 & n29185;
  assign n29187 = ~n11510 & n29186;
  assign n29188 = ~n10523 & n29187;
  assign n29189 = ~n11896 & n29188;
  assign n29190 = n11895 & n29189;
  assign n29191 = n11891 & n29190;
  assign n29192 = n11927 & n29191;
  assign n29193 = ~n29176 & ~n29192;
  assign n29194 = pi200 & ~n10939;
  assign n29195 = n12473 & n29194;
  assign n29196 = n12317 & n29195;
  assign n29197 = n12316 & n29196;
  assign n29198 = ~n11188 & n29197;
  assign n29199 = ~n12314 & n29198;
  assign n29200 = ~n11510 & n29199;
  assign n29201 = ~n11505 & n29200;
  assign n29202 = n11970 & n29201;
  assign n29203 = n12325 & n29202;
  assign n29204 = n12313 & n29203;
  assign n29205 = n12379 & n29204;
  assign n29206 = pi192 & ~n10074;
  assign n29207 = ~n11510 & n29206;
  assign n29208 = ~n11343 & n29207;
  assign n29209 = ~n11509 & n29208;
  assign n29210 = n11508 & n29209;
  assign n29211 = n11503 & n29210;
  assign n29212 = n11550 & n29211;
  assign n29213 = ~n29205 & ~n29212;
  assign n29214 = n29193 & n29213;
  assign n29215 = ~n9453 & n26982;
  assign n29216 = ~n11510 & n29215;
  assign n29217 = ~n10705 & n29216;
  assign n29218 = ~n12112 & n29217;
  assign n29219 = n12118 & n29218;
  assign n29220 = n11508 & n29219;
  assign n29221 = n12111 & n29220;
  assign n29222 = pi056 & ~n2176;
  assign n29223 = n4955 & n29222;
  assign n29224 = n7909 & n29223;
  assign n29225 = ~n2242 & n29224;
  assign n29226 = ~n3095 & n29225;
  assign n29227 = ~n3997 & n29226;
  assign n29228 = ~n4003 & n29227;
  assign n29229 = ~n4837 & n29228;
  assign n29230 = ~n5822 & n29229;
  assign n29231 = ~n6820 & n29230;
  assign n29232 = ~n7785 & n29231;
  assign n29233 = ~n9027 & n29232;
  assign n29234 = ~n10245 & n29233;
  assign n29235 = ~n11733 & n29234;
  assign n29236 = ~n11732 & n29235;
  assign n29237 = ~n11731 & n29236;
  assign n29238 = ~n11536 & n29237;
  assign n29239 = ~n11730 & n29238;
  assign n29240 = n11729 & n29239;
  assign n29241 = n11724 & n29240;
  assign n29242 = n11768 & n29241;
  assign n29243 = ~n29221 & ~n29242;
  assign n29244 = n12013 & n21872;
  assign n29245 = ~n5808 & n29244;
  assign n29246 = ~n6056 & n29245;
  assign n29247 = ~n7073 & n29246;
  assign n29248 = ~n8179 & n29247;
  assign n29249 = ~n9344 & n29248;
  assign n29250 = ~n11974 & n29249;
  assign n29251 = ~n11973 & n29250;
  assign n29252 = ~n11510 & n29251;
  assign n29253 = ~n10594 & n29252;
  assign n29254 = ~n11972 & n29253;
  assign n29255 = n11971 & n29254;
  assign n29256 = n11968 & n29255;
  assign n29257 = n12004 & n29256;
  assign n29258 = n12275 & n26923;
  assign n29259 = n11562 & n29258;
  assign n29260 = n11560 & n29259;
  assign n29261 = ~n9929 & n29260;
  assign n29262 = ~n11558 & n29261;
  assign n29263 = ~n11557 & n29262;
  assign n29264 = ~n11510 & n29263;
  assign n29265 = ~n11266 & n29264;
  assign n29266 = ~n11509 & n29265;
  assign n29267 = n11508 & n29266;
  assign n29268 = n11556 & n29267;
  assign n29269 = n11587 & n29268;
  assign n29270 = ~n29257 & ~n29269;
  assign n29271 = n29243 & n29270;
  assign n29272 = n29214 & n29271;
  assign n29273 = n29168 & n29272;
  assign po113 = ~n29116 | ~n29273;
  assign n29275 = ~n10460 & n27089;
  assign n29276 = ~n11510 & n29275;
  assign n29277 = ~n11852 & n29276;
  assign n29278 = n11859 & n29277;
  assign n29279 = ~n10400 & n27093;
  assign n29280 = ~n11790 & n29279;
  assign n29281 = n11795 & n29280;
  assign n29282 = pi225 & ~n501;
  assign n29283 = n12872 & n29282;
  assign n29284 = n14253 & n29283;
  assign n29285 = n12564 & n29284;
  assign n29286 = n28654 & n29285;
  assign n29287 = n12548 & n29286;
  assign n29288 = ~n1172 & n29287;
  assign n29289 = ~n996 & n29288;
  assign n29290 = ~n2306 & n29289;
  assign n29291 = n12571 & n29290;
  assign n29292 = n6677 & n29291;
  assign n29293 = n12580 & n29292;
  assign n29294 = n28668 & n29293;
  assign n29295 = n12542 & n29294;
  assign n29296 = n28650 & n29295;
  assign n29297 = ~n7236 & n29296;
  assign n29298 = ~n6137 & n29297;
  assign n29299 = n6193 & n29298;
  assign n29300 = n6134 & n29299;
  assign n29301 = ~n8867 & n29300;
  assign n29302 = ~n7235 & n29301;
  assign n29303 = n7296 & n29302;
  assign n29304 = n7231 & n29303;
  assign n29305 = ~n10027 & n29304;
  assign n29306 = ~n8866 & n29305;
  assign n29307 = n8898 & n29306;
  assign n29308 = n8863 & n29307;
  assign n29309 = pi217 & ~n501;
  assign n29310 = n12611 & n29309;
  assign n29311 = n26571 & n29310;
  assign n29312 = n12619 & n29311;
  assign n29313 = n28689 & n29312;
  assign n29314 = n12601 & n29313;
  assign n29315 = ~n1172 & n29314;
  assign n29316 = ~n996 & n29315;
  assign n29317 = ~n2306 & n29316;
  assign n29318 = n12626 & n29317;
  assign n29319 = n12628 & n29318;
  assign n29320 = n3823 & n29319;
  assign n29321 = n12634 & n29320;
  assign n29322 = n12682 & n29321;
  assign n29323 = n12844 & n29322;
  assign n29324 = ~n7236 & n29323;
  assign n29325 = ~n6137 & n29324;
  assign n29326 = n6193 & n29325;
  assign n29327 = n6134 & n29326;
  assign n29328 = ~n8867 & n29327;
  assign n29329 = ~n7235 & n29328;
  assign n29330 = n7296 & n29329;
  assign n29331 = n7231 & n29330;
  assign n29332 = ~n10027 & n29331;
  assign n29333 = ~n8866 & n29332;
  assign n29334 = n8898 & n29333;
  assign n29335 = n8863 & n29334;
  assign n29336 = ~n29308 & ~n29335;
  assign n29337 = ~n10788 & ~n29336;
  assign n29338 = ~n10026 & n29337;
  assign n29339 = n10072 & n29338;
  assign n29340 = n10021 & n29339;
  assign n29341 = ~n29281 & ~n29340;
  assign n29342 = ~n29278 & n29341;
  assign n29343 = ~n10554 & n27155;
  assign n29344 = ~n11510 & n29343;
  assign n29345 = ~n11506 & n29344;
  assign n29346 = n11957 & n29345;
  assign n29347 = n11952 & n29346;
  assign n29348 = ~n10629 & n27160;
  assign n29349 = ~n11510 & n29348;
  assign n29350 = n11970 & n29349;
  assign n29351 = n12039 & n29350;
  assign n29352 = n12034 & n29351;
  assign n29353 = ~n29347 & ~n29352;
  assign n29354 = n29342 & n29353;
  assign n29355 = ~n10094 & n27200;
  assign n29356 = ~n11510 & n29355;
  assign n29357 = ~n11318 & n29356;
  assign n29358 = ~n11501 & n29357;
  assign n29359 = n11508 & n29358;
  assign n29360 = n12175 & n29359;
  assign n29361 = n12168 & n29360;
  assign n29362 = pi057 & ~n2176;
  assign n29363 = n4955 & n29362;
  assign n29364 = n7909 & n29363;
  assign n29365 = ~n2242 & n29364;
  assign n29366 = ~n3095 & n29365;
  assign n29367 = ~n3997 & n29366;
  assign n29368 = ~n4003 & n29367;
  assign n29369 = ~n4837 & n29368;
  assign n29370 = ~n5822 & n29369;
  assign n29371 = ~n6820 & n29370;
  assign n29372 = ~n7785 & n29371;
  assign n29373 = ~n9027 & n29372;
  assign n29374 = ~n10245 & n29373;
  assign n29375 = ~n11733 & n29374;
  assign n29376 = ~n11732 & n29375;
  assign n29377 = ~n11731 & n29376;
  assign n29378 = ~n11536 & n29377;
  assign n29379 = ~n11730 & n29378;
  assign n29380 = n11729 & n29379;
  assign n29381 = n11724 & n29380;
  assign n29382 = n11768 & n29381;
  assign n29383 = ~n29361 & ~n29382;
  assign n29384 = n12275 & n27167;
  assign n29385 = n11562 & n29384;
  assign n29386 = n11560 & n29385;
  assign n29387 = ~n9929 & n29386;
  assign n29388 = ~n11558 & n29387;
  assign n29389 = ~n11557 & n29388;
  assign n29390 = ~n11510 & n29389;
  assign n29391 = ~n11266 & n29390;
  assign n29392 = ~n11509 & n29391;
  assign n29393 = n11508 & n29392;
  assign n29394 = n11556 & n29393;
  assign n29395 = n11587 & n29394;
  assign n29396 = n11681 & n27215;
  assign n29397 = n11680 & n29396;
  assign n29398 = ~n1372 & n29397;
  assign n29399 = ~n2243 & n29398;
  assign n29400 = ~n3104 & n29399;
  assign n29401 = ~n3971 & n29400;
  assign n29402 = ~n4003 & n29401;
  assign n29403 = ~n4872 & n29402;
  assign n29404 = ~n5801 & n29403;
  assign n29405 = ~n6739 & n29404;
  assign n29406 = ~n7807 & n29405;
  assign n29407 = ~n8989 & n29406;
  assign n29408 = ~n10273 & n29407;
  assign n29409 = ~n11678 & n29408;
  assign n29410 = ~n11677 & n29409;
  assign n29411 = ~n11676 & n29410;
  assign n29412 = ~n11499 & n29411;
  assign n29413 = ~n11675 & n29412;
  assign n29414 = n11674 & n29413;
  assign n29415 = n11669 & n29414;
  assign n29416 = n11716 & n29415;
  assign n29417 = ~n29395 & ~n29416;
  assign n29418 = n29383 & n29417;
  assign n29419 = n29354 & n29418;
  assign n29420 = n9115 & n22056;
  assign n29421 = ~n3066 & n29420;
  assign n29422 = ~n3983 & n29421;
  assign n29423 = ~n4003 & n29422;
  assign n29424 = ~n4024 & n29423;
  assign n29425 = ~n4999 & n29424;
  assign n29426 = ~n5827 & n29425;
  assign n29427 = ~n6893 & n29426;
  assign n29428 = ~n7890 & n29427;
  assign n29429 = ~n9131 & n29428;
  assign n29430 = ~n11627 & n29429;
  assign n29431 = ~n11626 & n29430;
  assign n29432 = ~n11625 & n29431;
  assign n29433 = ~n10278 & n29432;
  assign n29434 = ~n11624 & n29433;
  assign n29435 = n11623 & n29434;
  assign n29436 = n11618 & n29435;
  assign n29437 = n11661 & n29436;
  assign n29438 = n11378 & n25253;
  assign n29439 = n9942 & n29438;
  assign n29440 = ~n8834 & n29439;
  assign n29441 = ~n10002 & n29440;
  assign n29442 = ~n12212 & n29441;
  assign n29443 = ~n12211 & n29442;
  assign n29444 = ~n11510 & n29443;
  assign n29445 = ~n11297 & n29444;
  assign n29446 = ~n11478 & n29445;
  assign n29447 = n11508 & n29446;
  assign n29448 = n12210 & n29447;
  assign n29449 = n12239 & n29448;
  assign n29450 = ~n29437 & ~n29449;
  assign n29451 = n5085 & n27053;
  assign n29452 = n11931 & n29451;
  assign n29453 = ~n4817 & n29452;
  assign n29454 = ~n4902 & n29453;
  assign n29455 = ~n6001 & n29454;
  assign n29456 = ~n7014 & n29455;
  assign n29457 = ~n8114 & n29456;
  assign n29458 = ~n9276 & n29457;
  assign n29459 = ~n11898 & n29458;
  assign n29460 = ~n11897 & n29459;
  assign n29461 = ~n11510 & n29460;
  assign n29462 = ~n10523 & n29461;
  assign n29463 = ~n11896 & n29462;
  assign n29464 = n11895 & n29463;
  assign n29465 = n11891 & n29464;
  assign n29466 = n11927 & n29465;
  assign n29467 = pi201 & ~n10939;
  assign n29468 = n12473 & n29467;
  assign n29469 = n12317 & n29468;
  assign n29470 = n12316 & n29469;
  assign n29471 = ~n11188 & n29470;
  assign n29472 = ~n12314 & n29471;
  assign n29473 = ~n11510 & n29472;
  assign n29474 = ~n11505 & n29473;
  assign n29475 = n11970 & n29474;
  assign n29476 = n12325 & n29475;
  assign n29477 = n12313 & n29476;
  assign n29478 = n12379 & n29477;
  assign n29479 = ~n29466 & ~n29478;
  assign n29480 = n29450 & n29479;
  assign n29481 = ~n9533 & n27193;
  assign n29482 = ~n11510 & n29481;
  assign n29483 = ~n10787 & n29482;
  assign n29484 = ~n11478 & n29483;
  assign n29485 = n11593 & n29484;
  assign n29486 = n11508 & n29485;
  assign n29487 = n11610 & n29486;
  assign n29488 = n12182 & n23527;
  assign n29489 = ~n7869 & n29488;
  assign n29490 = ~n8346 & n29489;
  assign n29491 = ~n9485 & n29490;
  assign n29492 = ~n12130 & n29491;
  assign n29493 = ~n12129 & n29492;
  assign n29494 = ~n11510 & n29493;
  assign n29495 = ~n10741 & n29494;
  assign n29496 = ~n11501 & n29495;
  assign n29497 = n11508 & n29496;
  assign n29498 = n12128 & n29497;
  assign n29499 = n12157 & n29498;
  assign n29500 = ~n29487 & ~n29499;
  assign n29501 = n5062 & n27270;
  assign n29502 = n11861 & n29501;
  assign n29503 = ~n3940 & n29502;
  assign n29504 = ~n4001 & n29503;
  assign n29505 = ~n5043 & n29504;
  assign n29506 = ~n5943 & n29505;
  assign n29507 = ~n6951 & n29506;
  assign n29508 = ~n8037 & n29507;
  assign n29509 = ~n9200 & n29508;
  assign n29510 = ~n11813 & n29509;
  assign n29511 = ~n11812 & n29510;
  assign n29512 = ~n11510 & n29511;
  assign n29513 = ~n10445 & n29512;
  assign n29514 = ~n11811 & n29513;
  assign n29515 = n11810 & n29514;
  assign n29516 = n11805 & n29515;
  assign n29517 = n11845 & n29516;
  assign n29518 = pi193 & ~n10074;
  assign n29519 = ~n11510 & n29518;
  assign n29520 = ~n11343 & n29519;
  assign n29521 = ~n11509 & n29520;
  assign n29522 = n11508 & n29521;
  assign n29523 = n11503 & n29522;
  assign n29524 = n11550 & n29523;
  assign n29525 = ~n29517 & ~n29524;
  assign n29526 = n29500 & n29525;
  assign n29527 = pi209 & ~n10879;
  assign n29528 = ~n12412 & n29527;
  assign n29529 = ~n11510 & n29528;
  assign n29530 = ~n11505 & n29529;
  assign n29531 = n11970 & n29530;
  assign n29532 = n12325 & n29531;
  assign n29533 = n12411 & n29532;
  assign n29534 = n12470 & n29533;
  assign n29535 = n7177 & n27238;
  assign n29536 = n8261 & n29535;
  assign n29537 = ~n6784 & n29536;
  assign n29538 = ~n7158 & n29537;
  assign n29539 = ~n8250 & n29538;
  assign n29540 = ~n9414 & n29539;
  assign n29541 = ~n12053 & n29540;
  assign n29542 = ~n12052 & n29541;
  assign n29543 = ~n11510 & n29542;
  assign n29544 = ~n10667 & n29543;
  assign n29545 = ~n12051 & n29544;
  assign n29546 = n11508 & n29545;
  assign n29547 = n12050 & n29546;
  assign n29548 = n12082 & n29547;
  assign n29549 = ~n29534 & ~n29548;
  assign n29550 = ~n9453 & n27208;
  assign n29551 = ~n11510 & n29550;
  assign n29552 = ~n10705 & n29551;
  assign n29553 = ~n12112 & n29552;
  assign n29554 = n12118 & n29553;
  assign n29555 = n11508 & n29554;
  assign n29556 = n12111 & n29555;
  assign n29557 = n12013 & n22073;
  assign n29558 = ~n5808 & n29557;
  assign n29559 = ~n6056 & n29558;
  assign n29560 = ~n7073 & n29559;
  assign n29561 = ~n8179 & n29560;
  assign n29562 = ~n9344 & n29561;
  assign n29563 = ~n11974 & n29562;
  assign n29564 = ~n11973 & n29563;
  assign n29565 = ~n11510 & n29564;
  assign n29566 = ~n10594 & n29565;
  assign n29567 = ~n11972 & n29566;
  assign n29568 = n11971 & n29567;
  assign n29569 = n11968 & n29568;
  assign n29570 = n12004 & n29569;
  assign n29571 = ~n29556 & ~n29570;
  assign n29572 = n29549 & n29571;
  assign n29573 = n29526 & n29572;
  assign n29574 = n29480 & n29573;
  assign po114 = ~n29419 | ~n29574;
  assign n29576 = ~n10460 & n27357;
  assign n29577 = ~n11510 & n29576;
  assign n29578 = ~n11852 & n29577;
  assign n29579 = n11859 & n29578;
  assign n29580 = ~n10400 & n27361;
  assign n29581 = ~n11790 & n29580;
  assign n29582 = n11795 & n29581;
  assign n29583 = pi218 & ~n501;
  assign n29584 = n12611 & n29583;
  assign n29585 = n26571 & n29584;
  assign n29586 = n12619 & n29585;
  assign n29587 = n28689 & n29586;
  assign n29588 = n12601 & n29587;
  assign n29589 = ~n1172 & n29588;
  assign n29590 = ~n996 & n29589;
  assign n29591 = ~n2306 & n29590;
  assign n29592 = n12626 & n29591;
  assign n29593 = n12628 & n29592;
  assign n29594 = n3823 & n29593;
  assign n29595 = n12634 & n29594;
  assign n29596 = n12682 & n29595;
  assign n29597 = n12844 & n29596;
  assign n29598 = ~n7236 & n29597;
  assign n29599 = ~n6137 & n29598;
  assign n29600 = n6193 & n29599;
  assign n29601 = n6134 & n29600;
  assign n29602 = ~n8867 & n29601;
  assign n29603 = ~n7235 & n29602;
  assign n29604 = n7296 & n29603;
  assign n29605 = n7231 & n29604;
  assign n29606 = ~n10027 & n29605;
  assign n29607 = ~n8866 & n29606;
  assign n29608 = n8898 & n29607;
  assign n29609 = n8863 & n29608;
  assign n29610 = pi226 & ~n501;
  assign n29611 = n12872 & n29610;
  assign n29612 = n14253 & n29611;
  assign n29613 = n12564 & n29612;
  assign n29614 = n28654 & n29613;
  assign n29615 = n12548 & n29614;
  assign n29616 = ~n1172 & n29615;
  assign n29617 = ~n996 & n29616;
  assign n29618 = ~n2306 & n29617;
  assign n29619 = n12571 & n29618;
  assign n29620 = n6677 & n29619;
  assign n29621 = n12580 & n29620;
  assign n29622 = n28668 & n29621;
  assign n29623 = n12542 & n29622;
  assign n29624 = n28650 & n29623;
  assign n29625 = ~n7236 & n29624;
  assign n29626 = ~n6137 & n29625;
  assign n29627 = n6193 & n29626;
  assign n29628 = n6134 & n29627;
  assign n29629 = ~n8867 & n29628;
  assign n29630 = ~n7235 & n29629;
  assign n29631 = n7296 & n29630;
  assign n29632 = n7231 & n29631;
  assign n29633 = ~n10027 & n29632;
  assign n29634 = ~n8866 & n29633;
  assign n29635 = n8898 & n29634;
  assign n29636 = n8863 & n29635;
  assign n29637 = ~n29609 & ~n29636;
  assign n29638 = ~n10788 & ~n29637;
  assign n29639 = ~n10026 & n29638;
  assign n29640 = n10072 & n29639;
  assign n29641 = n10021 & n29640;
  assign n29642 = ~n29582 & ~n29641;
  assign n29643 = ~n29579 & n29642;
  assign n29644 = ~n10554 & n27423;
  assign n29645 = ~n11510 & n29644;
  assign n29646 = ~n11506 & n29645;
  assign n29647 = n11957 & n29646;
  assign n29648 = n11952 & n29647;
  assign n29649 = ~n10629 & n27428;
  assign n29650 = ~n11510 & n29649;
  assign n29651 = n11970 & n29650;
  assign n29652 = n12039 & n29651;
  assign n29653 = n12034 & n29652;
  assign n29654 = ~n29648 & ~n29653;
  assign n29655 = n29643 & n29654;
  assign n29656 = n12275 & n27344;
  assign n29657 = n11562 & n29656;
  assign n29658 = n11560 & n29657;
  assign n29659 = ~n9929 & n29658;
  assign n29660 = ~n11558 & n29659;
  assign n29661 = ~n11557 & n29660;
  assign n29662 = ~n11510 & n29661;
  assign n29663 = ~n11266 & n29662;
  assign n29664 = ~n11509 & n29663;
  assign n29665 = n11508 & n29664;
  assign n29666 = n11556 & n29665;
  assign n29667 = n11587 & n29666;
  assign n29668 = n11681 & n27477;
  assign n29669 = n11680 & n29668;
  assign n29670 = ~n1372 & n29669;
  assign n29671 = ~n2243 & n29670;
  assign n29672 = ~n3104 & n29671;
  assign n29673 = ~n3971 & n29672;
  assign n29674 = ~n4003 & n29673;
  assign n29675 = ~n4872 & n29674;
  assign n29676 = ~n5801 & n29675;
  assign n29677 = ~n6739 & n29676;
  assign n29678 = ~n7807 & n29677;
  assign n29679 = ~n8989 & n29678;
  assign n29680 = ~n10273 & n29679;
  assign n29681 = ~n11678 & n29680;
  assign n29682 = ~n11677 & n29681;
  assign n29683 = ~n11676 & n29682;
  assign n29684 = ~n11499 & n29683;
  assign n29685 = ~n11675 & n29684;
  assign n29686 = n11674 & n29685;
  assign n29687 = n11669 & n29686;
  assign n29688 = n11716 & n29687;
  assign n29689 = ~n29667 & ~n29688;
  assign n29690 = pi058 & ~n2176;
  assign n29691 = n4955 & n29690;
  assign n29692 = n7909 & n29691;
  assign n29693 = ~n2242 & n29692;
  assign n29694 = ~n3095 & n29693;
  assign n29695 = ~n3997 & n29694;
  assign n29696 = ~n4003 & n29695;
  assign n29697 = ~n4837 & n29696;
  assign n29698 = ~n5822 & n29697;
  assign n29699 = ~n6820 & n29698;
  assign n29700 = ~n7785 & n29699;
  assign n29701 = ~n9027 & n29700;
  assign n29702 = ~n10245 & n29701;
  assign n29703 = ~n11733 & n29702;
  assign n29704 = ~n11732 & n29703;
  assign n29705 = ~n11731 & n29704;
  assign n29706 = ~n11536 & n29705;
  assign n29707 = ~n11730 & n29706;
  assign n29708 = n11729 & n29707;
  assign n29709 = n11724 & n29708;
  assign n29710 = n11768 & n29709;
  assign n29711 = ~n9453 & n27470;
  assign n29712 = ~n11510 & n29711;
  assign n29713 = ~n10705 & n29712;
  assign n29714 = ~n12112 & n29713;
  assign n29715 = n12118 & n29714;
  assign n29716 = n11508 & n29715;
  assign n29717 = n12111 & n29716;
  assign n29718 = ~n29710 & ~n29717;
  assign n29719 = n29689 & n29718;
  assign n29720 = n29655 & n29719;
  assign n29721 = n9115 & n22281;
  assign n29722 = ~n3066 & n29721;
  assign n29723 = ~n3983 & n29722;
  assign n29724 = ~n4003 & n29723;
  assign n29725 = ~n4024 & n29724;
  assign n29726 = ~n4999 & n29725;
  assign n29727 = ~n5827 & n29726;
  assign n29728 = ~n6893 & n29727;
  assign n29729 = ~n7890 & n29728;
  assign n29730 = ~n9131 & n29729;
  assign n29731 = ~n11627 & n29730;
  assign n29732 = ~n11626 & n29731;
  assign n29733 = ~n11625 & n29732;
  assign n29734 = ~n10278 & n29733;
  assign n29735 = ~n11624 & n29734;
  assign n29736 = n11623 & n29735;
  assign n29737 = n11618 & n29736;
  assign n29738 = n11661 & n29737;
  assign n29739 = n11378 & n25513;
  assign n29740 = n9942 & n29739;
  assign n29741 = ~n8834 & n29740;
  assign n29742 = ~n10002 & n29741;
  assign n29743 = ~n12212 & n29742;
  assign n29744 = ~n12211 & n29743;
  assign n29745 = ~n11510 & n29744;
  assign n29746 = ~n11297 & n29745;
  assign n29747 = ~n11478 & n29746;
  assign n29748 = n11508 & n29747;
  assign n29749 = n12210 & n29748;
  assign n29750 = n12239 & n29749;
  assign n29751 = ~n29738 & ~n29750;
  assign n29752 = n5085 & n27537;
  assign n29753 = n11931 & n29752;
  assign n29754 = ~n4817 & n29753;
  assign n29755 = ~n4902 & n29754;
  assign n29756 = ~n6001 & n29755;
  assign n29757 = ~n7014 & n29756;
  assign n29758 = ~n8114 & n29757;
  assign n29759 = ~n9276 & n29758;
  assign n29760 = ~n11898 & n29759;
  assign n29761 = ~n11897 & n29760;
  assign n29762 = ~n11510 & n29761;
  assign n29763 = ~n10523 & n29762;
  assign n29764 = ~n11896 & n29763;
  assign n29765 = n11895 & n29764;
  assign n29766 = n11891 & n29765;
  assign n29767 = n11927 & n29766;
  assign n29768 = pi202 & ~n10939;
  assign n29769 = n12473 & n29768;
  assign n29770 = n12317 & n29769;
  assign n29771 = n12316 & n29770;
  assign n29772 = ~n11188 & n29771;
  assign n29773 = ~n12314 & n29772;
  assign n29774 = ~n11510 & n29773;
  assign n29775 = ~n11505 & n29774;
  assign n29776 = n11970 & n29775;
  assign n29777 = n12325 & n29776;
  assign n29778 = n12313 & n29777;
  assign n29779 = n12379 & n29778;
  assign n29780 = ~n29767 & ~n29779;
  assign n29781 = n29751 & n29780;
  assign n29782 = ~n10094 & n27337;
  assign n29783 = ~n11510 & n29782;
  assign n29784 = ~n11318 & n29783;
  assign n29785 = ~n11501 & n29784;
  assign n29786 = n11508 & n29785;
  assign n29787 = n12175 & n29786;
  assign n29788 = n12168 & n29787;
  assign n29789 = n12182 & n23753;
  assign n29790 = ~n7869 & n29789;
  assign n29791 = ~n8346 & n29790;
  assign n29792 = ~n9485 & n29791;
  assign n29793 = ~n12130 & n29792;
  assign n29794 = ~n12129 & n29793;
  assign n29795 = ~n11510 & n29794;
  assign n29796 = ~n10741 & n29795;
  assign n29797 = ~n11501 & n29796;
  assign n29798 = n11508 & n29797;
  assign n29799 = n12128 & n29798;
  assign n29800 = n12157 & n29799;
  assign n29801 = ~n29788 & ~n29800;
  assign n29802 = pi194 & ~n10074;
  assign n29803 = ~n11510 & n29802;
  assign n29804 = ~n11343 & n29803;
  assign n29805 = ~n11509 & n29804;
  assign n29806 = n11508 & n29805;
  assign n29807 = n11503 & n29806;
  assign n29808 = n11550 & n29807;
  assign n29809 = n5062 & n27506;
  assign n29810 = n11861 & n29809;
  assign n29811 = ~n3940 & n29810;
  assign n29812 = ~n4001 & n29811;
  assign n29813 = ~n5043 & n29812;
  assign n29814 = ~n5943 & n29813;
  assign n29815 = ~n6951 & n29814;
  assign n29816 = ~n8037 & n29815;
  assign n29817 = ~n9200 & n29816;
  assign n29818 = ~n11813 & n29817;
  assign n29819 = ~n11812 & n29818;
  assign n29820 = ~n11510 & n29819;
  assign n29821 = ~n10445 & n29820;
  assign n29822 = ~n11811 & n29821;
  assign n29823 = n11810 & n29822;
  assign n29824 = n11805 & n29823;
  assign n29825 = n11845 & n29824;
  assign n29826 = ~n29808 & ~n29825;
  assign n29827 = n29801 & n29826;
  assign n29828 = ~n9533 & n27499;
  assign n29829 = ~n11510 & n29828;
  assign n29830 = ~n10787 & n29829;
  assign n29831 = ~n11478 & n29830;
  assign n29832 = n11593 & n29831;
  assign n29833 = n11508 & n29832;
  assign n29834 = n11610 & n29833;
  assign n29835 = n7177 & n27435;
  assign n29836 = n8261 & n29835;
  assign n29837 = ~n6784 & n29836;
  assign n29838 = ~n7158 & n29837;
  assign n29839 = ~n8250 & n29838;
  assign n29840 = ~n9414 & n29839;
  assign n29841 = ~n12053 & n29840;
  assign n29842 = ~n12052 & n29841;
  assign n29843 = ~n11510 & n29842;
  assign n29844 = ~n10667 & n29843;
  assign n29845 = ~n12051 & n29844;
  assign n29846 = n11508 & n29845;
  assign n29847 = n12050 & n29846;
  assign n29848 = n12082 & n29847;
  assign n29849 = ~n29834 & ~n29848;
  assign n29850 = n12013 & n22231;
  assign n29851 = ~n5808 & n29850;
  assign n29852 = ~n6056 & n29851;
  assign n29853 = ~n7073 & n29852;
  assign n29854 = ~n8179 & n29853;
  assign n29855 = ~n9344 & n29854;
  assign n29856 = ~n11974 & n29855;
  assign n29857 = ~n11973 & n29856;
  assign n29858 = ~n11510 & n29857;
  assign n29859 = ~n10594 & n29858;
  assign n29860 = ~n11972 & n29859;
  assign n29861 = n11971 & n29860;
  assign n29862 = n11968 & n29861;
  assign n29863 = n12004 & n29862;
  assign n29864 = pi210 & ~n10879;
  assign n29865 = ~n12412 & n29864;
  assign n29866 = ~n11510 & n29865;
  assign n29867 = ~n11505 & n29866;
  assign n29868 = n11970 & n29867;
  assign n29869 = n12325 & n29868;
  assign n29870 = n12411 & n29869;
  assign n29871 = n12470 & n29870;
  assign n29872 = ~n29863 & ~n29871;
  assign n29873 = n29849 & n29872;
  assign n29874 = n29827 & n29873;
  assign n29875 = n29781 & n29874;
  assign po115 = ~n29720 | ~n29875;
  assign n29877 = ~n10460 & n27621;
  assign n29878 = ~n11510 & n29877;
  assign n29879 = ~n11852 & n29878;
  assign n29880 = n11859 & n29879;
  assign n29881 = ~n10400 & n27625;
  assign n29882 = ~n11790 & n29881;
  assign n29883 = n11795 & n29882;
  assign n29884 = pi227 & ~n501;
  assign n29885 = n12872 & n29884;
  assign n29886 = n14253 & n29885;
  assign n29887 = n12564 & n29886;
  assign n29888 = n28654 & n29887;
  assign n29889 = n12548 & n29888;
  assign n29890 = ~n1172 & n29889;
  assign n29891 = ~n996 & n29890;
  assign n29892 = ~n2306 & n29891;
  assign n29893 = n12571 & n29892;
  assign n29894 = n6677 & n29893;
  assign n29895 = n12580 & n29894;
  assign n29896 = n28668 & n29895;
  assign n29897 = n12542 & n29896;
  assign n29898 = n28650 & n29897;
  assign n29899 = ~n7236 & n29898;
  assign n29900 = ~n6137 & n29899;
  assign n29901 = n6193 & n29900;
  assign n29902 = n6134 & n29901;
  assign n29903 = ~n8867 & n29902;
  assign n29904 = ~n7235 & n29903;
  assign n29905 = n7296 & n29904;
  assign n29906 = n7231 & n29905;
  assign n29907 = ~n10027 & n29906;
  assign n29908 = ~n8866 & n29907;
  assign n29909 = n8898 & n29908;
  assign n29910 = n8863 & n29909;
  assign n29911 = pi219 & ~n501;
  assign n29912 = n12611 & n29911;
  assign n29913 = n26571 & n29912;
  assign n29914 = n12619 & n29913;
  assign n29915 = n28689 & n29914;
  assign n29916 = n12601 & n29915;
  assign n29917 = ~n1172 & n29916;
  assign n29918 = ~n996 & n29917;
  assign n29919 = ~n2306 & n29918;
  assign n29920 = n12626 & n29919;
  assign n29921 = n12628 & n29920;
  assign n29922 = n3823 & n29921;
  assign n29923 = n12634 & n29922;
  assign n29924 = n12682 & n29923;
  assign n29925 = n12844 & n29924;
  assign n29926 = ~n7236 & n29925;
  assign n29927 = ~n6137 & n29926;
  assign n29928 = n6193 & n29927;
  assign n29929 = n6134 & n29928;
  assign n29930 = ~n8867 & n29929;
  assign n29931 = ~n7235 & n29930;
  assign n29932 = n7296 & n29931;
  assign n29933 = n7231 & n29932;
  assign n29934 = ~n10027 & n29933;
  assign n29935 = ~n8866 & n29934;
  assign n29936 = n8898 & n29935;
  assign n29937 = n8863 & n29936;
  assign n29938 = ~n29910 & ~n29937;
  assign n29939 = ~n10788 & ~n29938;
  assign n29940 = ~n10026 & n29939;
  assign n29941 = n10072 & n29940;
  assign n29942 = n10021 & n29941;
  assign n29943 = ~n29883 & ~n29942;
  assign n29944 = ~n29880 & n29943;
  assign n29945 = ~n10554 & n27687;
  assign n29946 = ~n11510 & n29945;
  assign n29947 = ~n11506 & n29946;
  assign n29948 = n11957 & n29947;
  assign n29949 = n11952 & n29948;
  assign n29950 = ~n10629 & n27692;
  assign n29951 = ~n11510 & n29950;
  assign n29952 = n11970 & n29951;
  assign n29953 = n12039 & n29952;
  assign n29954 = n12034 & n29953;
  assign n29955 = ~n29949 & ~n29954;
  assign n29956 = n29944 & n29955;
  assign n29957 = n12275 & n27608;
  assign n29958 = n11562 & n29957;
  assign n29959 = n11560 & n29958;
  assign n29960 = ~n9929 & n29959;
  assign n29961 = ~n11558 & n29960;
  assign n29962 = ~n11557 & n29961;
  assign n29963 = ~n11510 & n29962;
  assign n29964 = ~n11266 & n29963;
  assign n29965 = ~n11509 & n29964;
  assign n29966 = n11508 & n29965;
  assign n29967 = n11556 & n29966;
  assign n29968 = n11587 & n29967;
  assign n29969 = n11681 & n27731;
  assign n29970 = n11680 & n29969;
  assign n29971 = ~n1372 & n29970;
  assign n29972 = ~n2243 & n29971;
  assign n29973 = ~n3104 & n29972;
  assign n29974 = ~n3971 & n29973;
  assign n29975 = ~n4003 & n29974;
  assign n29976 = ~n4872 & n29975;
  assign n29977 = ~n5801 & n29976;
  assign n29978 = ~n6739 & n29977;
  assign n29979 = ~n7807 & n29978;
  assign n29980 = ~n8989 & n29979;
  assign n29981 = ~n10273 & n29980;
  assign n29982 = ~n11678 & n29981;
  assign n29983 = ~n11677 & n29982;
  assign n29984 = ~n11676 & n29983;
  assign n29985 = ~n11499 & n29984;
  assign n29986 = ~n11675 & n29985;
  assign n29987 = n11674 & n29986;
  assign n29988 = n11669 & n29987;
  assign n29989 = n11716 & n29988;
  assign n29990 = ~n29968 & ~n29989;
  assign n29991 = pi059 & ~n2176;
  assign n29992 = n4955 & n29991;
  assign n29993 = n7909 & n29992;
  assign n29994 = ~n2242 & n29993;
  assign n29995 = ~n3095 & n29994;
  assign n29996 = ~n3997 & n29995;
  assign n29997 = ~n4003 & n29996;
  assign n29998 = ~n4837 & n29997;
  assign n29999 = ~n5822 & n29998;
  assign n30000 = ~n6820 & n29999;
  assign n30001 = ~n7785 & n30000;
  assign n30002 = ~n9027 & n30001;
  assign n30003 = ~n10245 & n30002;
  assign n30004 = ~n11733 & n30003;
  assign n30005 = ~n11732 & n30004;
  assign n30006 = ~n11731 & n30005;
  assign n30007 = ~n11536 & n30006;
  assign n30008 = ~n11730 & n30007;
  assign n30009 = n11729 & n30008;
  assign n30010 = n11724 & n30009;
  assign n30011 = n11768 & n30010;
  assign n30012 = n12013 & n22398;
  assign n30013 = ~n5808 & n30012;
  assign n30014 = ~n6056 & n30013;
  assign n30015 = ~n7073 & n30014;
  assign n30016 = ~n8179 & n30015;
  assign n30017 = ~n9344 & n30016;
  assign n30018 = ~n11974 & n30017;
  assign n30019 = ~n11973 & n30018;
  assign n30020 = ~n11510 & n30019;
  assign n30021 = ~n10594 & n30020;
  assign n30022 = ~n11972 & n30021;
  assign n30023 = n11971 & n30022;
  assign n30024 = n11968 & n30023;
  assign n30025 = n12004 & n30024;
  assign n30026 = ~n30011 & ~n30025;
  assign n30027 = n29990 & n30026;
  assign n30028 = n29956 & n30027;
  assign n30029 = n5085 & n27803;
  assign n30030 = n11931 & n30029;
  assign n30031 = ~n4817 & n30030;
  assign n30032 = ~n4902 & n30031;
  assign n30033 = ~n6001 & n30032;
  assign n30034 = ~n7014 & n30033;
  assign n30035 = ~n8114 & n30034;
  assign n30036 = ~n9276 & n30035;
  assign n30037 = ~n11898 & n30036;
  assign n30038 = ~n11897 & n30037;
  assign n30039 = ~n11510 & n30038;
  assign n30040 = ~n10523 & n30039;
  assign n30041 = ~n11896 & n30040;
  assign n30042 = n11895 & n30041;
  assign n30043 = n11891 & n30042;
  assign n30044 = n11927 & n30043;
  assign n30045 = n11378 & n25600;
  assign n30046 = n9942 & n30045;
  assign n30047 = ~n8834 & n30046;
  assign n30048 = ~n10002 & n30047;
  assign n30049 = ~n12212 & n30048;
  assign n30050 = ~n12211 & n30049;
  assign n30051 = ~n11510 & n30050;
  assign n30052 = ~n11297 & n30051;
  assign n30053 = ~n11478 & n30052;
  assign n30054 = n11508 & n30053;
  assign n30055 = n12210 & n30054;
  assign n30056 = n12239 & n30055;
  assign n30057 = ~n30044 & ~n30056;
  assign n30058 = n9115 & n22448;
  assign n30059 = ~n3066 & n30058;
  assign n30060 = ~n3983 & n30059;
  assign n30061 = ~n4003 & n30060;
  assign n30062 = ~n4024 & n30061;
  assign n30063 = ~n4999 & n30062;
  assign n30064 = ~n5827 & n30063;
  assign n30065 = ~n6893 & n30064;
  assign n30066 = ~n7890 & n30065;
  assign n30067 = ~n9131 & n30066;
  assign n30068 = ~n11627 & n30067;
  assign n30069 = ~n11626 & n30068;
  assign n30070 = ~n11625 & n30069;
  assign n30071 = ~n10278 & n30070;
  assign n30072 = ~n11624 & n30071;
  assign n30073 = n11623 & n30072;
  assign n30074 = n11618 & n30073;
  assign n30075 = n11661 & n30074;
  assign n30076 = pi195 & ~n10074;
  assign n30077 = ~n11510 & n30076;
  assign n30078 = ~n11343 & n30077;
  assign n30079 = ~n11509 & n30078;
  assign n30080 = n11508 & n30079;
  assign n30081 = n11503 & n30080;
  assign n30082 = n11550 & n30081;
  assign n30083 = ~n30075 & ~n30082;
  assign n30084 = n30057 & n30083;
  assign n30085 = pi211 & ~n10879;
  assign n30086 = ~n12412 & n30085;
  assign n30087 = ~n11510 & n30086;
  assign n30088 = ~n11505 & n30087;
  assign n30089 = n11970 & n30088;
  assign n30090 = n12325 & n30089;
  assign n30091 = n12411 & n30090;
  assign n30092 = n12470 & n30091;
  assign n30093 = n12182 & n23946;
  assign n30094 = ~n7869 & n30093;
  assign n30095 = ~n8346 & n30094;
  assign n30096 = ~n9485 & n30095;
  assign n30097 = ~n12130 & n30096;
  assign n30098 = ~n12129 & n30097;
  assign n30099 = ~n11510 & n30098;
  assign n30100 = ~n10741 & n30099;
  assign n30101 = ~n11501 & n30100;
  assign n30102 = n11508 & n30101;
  assign n30103 = n12128 & n30102;
  assign n30104 = n12157 & n30103;
  assign n30105 = ~n30092 & ~n30104;
  assign n30106 = pi203 & ~n10939;
  assign n30107 = n12473 & n30106;
  assign n30108 = n12317 & n30107;
  assign n30109 = n12316 & n30108;
  assign n30110 = ~n11188 & n30109;
  assign n30111 = ~n12314 & n30110;
  assign n30112 = ~n11510 & n30111;
  assign n30113 = ~n11505 & n30112;
  assign n30114 = n11970 & n30113;
  assign n30115 = n12325 & n30114;
  assign n30116 = n12313 & n30115;
  assign n30117 = n12379 & n30116;
  assign n30118 = n5062 & n27770;
  assign n30119 = n11861 & n30118;
  assign n30120 = ~n3940 & n30119;
  assign n30121 = ~n4001 & n30120;
  assign n30122 = ~n5043 & n30121;
  assign n30123 = ~n5943 & n30122;
  assign n30124 = ~n6951 & n30123;
  assign n30125 = ~n8037 & n30124;
  assign n30126 = ~n9200 & n30125;
  assign n30127 = ~n11813 & n30126;
  assign n30128 = ~n11812 & n30127;
  assign n30129 = ~n11510 & n30128;
  assign n30130 = ~n10445 & n30129;
  assign n30131 = ~n11811 & n30130;
  assign n30132 = n11810 & n30131;
  assign n30133 = n11805 & n30132;
  assign n30134 = n11845 & n30133;
  assign n30135 = ~n30117 & ~n30134;
  assign n30136 = n30105 & n30135;
  assign n30137 = ~n9533 & n27593;
  assign n30138 = ~n11510 & n30137;
  assign n30139 = ~n10787 & n30138;
  assign n30140 = ~n11478 & n30139;
  assign n30141 = n11593 & n30140;
  assign n30142 = n11508 & n30141;
  assign n30143 = n11610 & n30142;
  assign n30144 = n7177 & n27789;
  assign n30145 = n8261 & n30144;
  assign n30146 = ~n6784 & n30145;
  assign n30147 = ~n7158 & n30146;
  assign n30148 = ~n8250 & n30147;
  assign n30149 = ~n9414 & n30148;
  assign n30150 = ~n12053 & n30149;
  assign n30151 = ~n12052 & n30150;
  assign n30152 = ~n11510 & n30151;
  assign n30153 = ~n10667 & n30152;
  assign n30154 = ~n12051 & n30153;
  assign n30155 = n11508 & n30154;
  assign n30156 = n12050 & n30155;
  assign n30157 = n12082 & n30156;
  assign n30158 = ~n30143 & ~n30157;
  assign n30159 = ~n10094 & n27601;
  assign n30160 = ~n11510 & n30159;
  assign n30161 = ~n11318 & n30160;
  assign n30162 = ~n11501 & n30161;
  assign n30163 = n11508 & n30162;
  assign n30164 = n12175 & n30163;
  assign n30165 = n12168 & n30164;
  assign n30166 = ~n9453 & n27724;
  assign n30167 = ~n11510 & n30166;
  assign n30168 = ~n10705 & n30167;
  assign n30169 = ~n12112 & n30168;
  assign n30170 = n12118 & n30169;
  assign n30171 = n11508 & n30170;
  assign n30172 = n12111 & n30171;
  assign n30173 = ~n30165 & ~n30172;
  assign n30174 = n30158 & n30173;
  assign n30175 = n30136 & n30174;
  assign n30176 = n30084 & n30175;
  assign po116 = ~n30028 | ~n30176;
  assign n30178 = ~n10460 & n27887;
  assign n30179 = ~n11510 & n30178;
  assign n30180 = ~n11852 & n30179;
  assign n30181 = n11859 & n30180;
  assign n30182 = ~n10400 & n27891;
  assign n30183 = ~n11790 & n30182;
  assign n30184 = n11795 & n30183;
  assign n30185 = pi228 & ~n501;
  assign n30186 = n12872 & n30185;
  assign n30187 = n14253 & n30186;
  assign n30188 = n12564 & n30187;
  assign n30189 = n28654 & n30188;
  assign n30190 = n12548 & n30189;
  assign n30191 = ~n1172 & n30190;
  assign n30192 = ~n996 & n30191;
  assign n30193 = ~n2306 & n30192;
  assign n30194 = n12571 & n30193;
  assign n30195 = n6677 & n30194;
  assign n30196 = n12580 & n30195;
  assign n30197 = n28668 & n30196;
  assign n30198 = n12542 & n30197;
  assign n30199 = n28650 & n30198;
  assign n30200 = ~n7236 & n30199;
  assign n30201 = ~n6137 & n30200;
  assign n30202 = n6193 & n30201;
  assign n30203 = n6134 & n30202;
  assign n30204 = ~n8867 & n30203;
  assign n30205 = ~n7235 & n30204;
  assign n30206 = n7296 & n30205;
  assign n30207 = n7231 & n30206;
  assign n30208 = ~n10027 & n30207;
  assign n30209 = ~n8866 & n30208;
  assign n30210 = n8898 & n30209;
  assign n30211 = n8863 & n30210;
  assign n30212 = pi220 & ~n501;
  assign n30213 = n12611 & n30212;
  assign n30214 = n26571 & n30213;
  assign n30215 = n12619 & n30214;
  assign n30216 = n28689 & n30215;
  assign n30217 = n12601 & n30216;
  assign n30218 = ~n1172 & n30217;
  assign n30219 = ~n996 & n30218;
  assign n30220 = ~n2306 & n30219;
  assign n30221 = n12626 & n30220;
  assign n30222 = n12628 & n30221;
  assign n30223 = n3823 & n30222;
  assign n30224 = n12634 & n30223;
  assign n30225 = n12682 & n30224;
  assign n30226 = n12844 & n30225;
  assign n30227 = ~n7236 & n30226;
  assign n30228 = ~n6137 & n30227;
  assign n30229 = n6193 & n30228;
  assign n30230 = n6134 & n30229;
  assign n30231 = ~n8867 & n30230;
  assign n30232 = ~n7235 & n30231;
  assign n30233 = n7296 & n30232;
  assign n30234 = n7231 & n30233;
  assign n30235 = ~n10027 & n30234;
  assign n30236 = ~n8866 & n30235;
  assign n30237 = n8898 & n30236;
  assign n30238 = n8863 & n30237;
  assign n30239 = ~n30211 & ~n30238;
  assign n30240 = ~n10788 & ~n30239;
  assign n30241 = ~n10026 & n30240;
  assign n30242 = n10072 & n30241;
  assign n30243 = n10021 & n30242;
  assign n30244 = ~n30184 & ~n30243;
  assign n30245 = ~n30181 & n30244;
  assign n30246 = ~n10554 & n27953;
  assign n30247 = ~n11510 & n30246;
  assign n30248 = ~n11506 & n30247;
  assign n30249 = n11957 & n30248;
  assign n30250 = n11952 & n30249;
  assign n30251 = ~n10629 & n27958;
  assign n30252 = ~n11510 & n30251;
  assign n30253 = n11970 & n30252;
  assign n30254 = n12039 & n30253;
  assign n30255 = n12034 & n30254;
  assign n30256 = ~n30250 & ~n30255;
  assign n30257 = n30245 & n30256;
  assign n30258 = n12275 & n27874;
  assign n30259 = n11562 & n30258;
  assign n30260 = n11560 & n30259;
  assign n30261 = ~n9929 & n30260;
  assign n30262 = ~n11558 & n30261;
  assign n30263 = ~n11557 & n30262;
  assign n30264 = ~n11510 & n30263;
  assign n30265 = ~n11266 & n30264;
  assign n30266 = ~n11509 & n30265;
  assign n30267 = n11508 & n30266;
  assign n30268 = n11556 & n30267;
  assign n30269 = n11587 & n30268;
  assign n30270 = n11681 & n27997;
  assign n30271 = n11680 & n30270;
  assign n30272 = ~n1372 & n30271;
  assign n30273 = ~n2243 & n30272;
  assign n30274 = ~n3104 & n30273;
  assign n30275 = ~n3971 & n30274;
  assign n30276 = ~n4003 & n30275;
  assign n30277 = ~n4872 & n30276;
  assign n30278 = ~n5801 & n30277;
  assign n30279 = ~n6739 & n30278;
  assign n30280 = ~n7807 & n30279;
  assign n30281 = ~n8989 & n30280;
  assign n30282 = ~n10273 & n30281;
  assign n30283 = ~n11678 & n30282;
  assign n30284 = ~n11677 & n30283;
  assign n30285 = ~n11676 & n30284;
  assign n30286 = ~n11499 & n30285;
  assign n30287 = ~n11675 & n30286;
  assign n30288 = n11674 & n30287;
  assign n30289 = n11669 & n30288;
  assign n30290 = n11716 & n30289;
  assign n30291 = ~n30269 & ~n30290;
  assign n30292 = pi060 & ~n2176;
  assign n30293 = n4955 & n30292;
  assign n30294 = n7909 & n30293;
  assign n30295 = ~n2242 & n30294;
  assign n30296 = ~n3095 & n30295;
  assign n30297 = ~n3997 & n30296;
  assign n30298 = ~n4003 & n30297;
  assign n30299 = ~n4837 & n30298;
  assign n30300 = ~n5822 & n30299;
  assign n30301 = ~n6820 & n30300;
  assign n30302 = ~n7785 & n30301;
  assign n30303 = ~n9027 & n30302;
  assign n30304 = ~n10245 & n30303;
  assign n30305 = ~n11733 & n30304;
  assign n30306 = ~n11732 & n30305;
  assign n30307 = ~n11731 & n30306;
  assign n30308 = ~n11536 & n30307;
  assign n30309 = ~n11730 & n30308;
  assign n30310 = n11729 & n30309;
  assign n30311 = n11724 & n30310;
  assign n30312 = n11768 & n30311;
  assign n30313 = n12013 & n22565;
  assign n30314 = ~n5808 & n30313;
  assign n30315 = ~n6056 & n30314;
  assign n30316 = ~n7073 & n30315;
  assign n30317 = ~n8179 & n30316;
  assign n30318 = ~n9344 & n30317;
  assign n30319 = ~n11974 & n30318;
  assign n30320 = ~n11973 & n30319;
  assign n30321 = ~n11510 & n30320;
  assign n30322 = ~n10594 & n30321;
  assign n30323 = ~n11972 & n30322;
  assign n30324 = n11971 & n30323;
  assign n30325 = n11968 & n30324;
  assign n30326 = n12004 & n30325;
  assign n30327 = ~n30312 & ~n30326;
  assign n30328 = n30291 & n30327;
  assign n30329 = n30257 & n30328;
  assign n30330 = n5085 & n28069;
  assign n30331 = n11931 & n30330;
  assign n30332 = ~n4817 & n30331;
  assign n30333 = ~n4902 & n30332;
  assign n30334 = ~n6001 & n30333;
  assign n30335 = ~n7014 & n30334;
  assign n30336 = ~n8114 & n30335;
  assign n30337 = ~n9276 & n30336;
  assign n30338 = ~n11898 & n30337;
  assign n30339 = ~n11897 & n30338;
  assign n30340 = ~n11510 & n30339;
  assign n30341 = ~n10523 & n30340;
  assign n30342 = ~n11896 & n30341;
  assign n30343 = n11895 & n30342;
  assign n30344 = n11891 & n30343;
  assign n30345 = n11927 & n30344;
  assign n30346 = n11378 & n25833;
  assign n30347 = n9942 & n30346;
  assign n30348 = ~n8834 & n30347;
  assign n30349 = ~n10002 & n30348;
  assign n30350 = ~n12212 & n30349;
  assign n30351 = ~n12211 & n30350;
  assign n30352 = ~n11510 & n30351;
  assign n30353 = ~n11297 & n30352;
  assign n30354 = ~n11478 & n30353;
  assign n30355 = n11508 & n30354;
  assign n30356 = n12210 & n30355;
  assign n30357 = n12239 & n30356;
  assign n30358 = ~n30345 & ~n30357;
  assign n30359 = n9115 & n22615;
  assign n30360 = ~n3066 & n30359;
  assign n30361 = ~n3983 & n30360;
  assign n30362 = ~n4003 & n30361;
  assign n30363 = ~n4024 & n30362;
  assign n30364 = ~n4999 & n30363;
  assign n30365 = ~n5827 & n30364;
  assign n30366 = ~n6893 & n30365;
  assign n30367 = ~n7890 & n30366;
  assign n30368 = ~n9131 & n30367;
  assign n30369 = ~n11627 & n30368;
  assign n30370 = ~n11626 & n30369;
  assign n30371 = ~n11625 & n30370;
  assign n30372 = ~n10278 & n30371;
  assign n30373 = ~n11624 & n30372;
  assign n30374 = n11623 & n30373;
  assign n30375 = n11618 & n30374;
  assign n30376 = n11661 & n30375;
  assign n30377 = pi196 & ~n10074;
  assign n30378 = ~n11510 & n30377;
  assign n30379 = ~n11343 & n30378;
  assign n30380 = ~n11509 & n30379;
  assign n30381 = n11508 & n30380;
  assign n30382 = n11503 & n30381;
  assign n30383 = n11550 & n30382;
  assign n30384 = ~n30376 & ~n30383;
  assign n30385 = n30358 & n30384;
  assign n30386 = pi212 & ~n10879;
  assign n30387 = ~n12412 & n30386;
  assign n30388 = ~n11510 & n30387;
  assign n30389 = ~n11505 & n30388;
  assign n30390 = n11970 & n30389;
  assign n30391 = n12325 & n30390;
  assign n30392 = n12411 & n30391;
  assign n30393 = n12470 & n30392;
  assign n30394 = n12182 & n24207;
  assign n30395 = ~n7869 & n30394;
  assign n30396 = ~n8346 & n30395;
  assign n30397 = ~n9485 & n30396;
  assign n30398 = ~n12130 & n30397;
  assign n30399 = ~n12129 & n30398;
  assign n30400 = ~n11510 & n30399;
  assign n30401 = ~n10741 & n30400;
  assign n30402 = ~n11501 & n30401;
  assign n30403 = n11508 & n30402;
  assign n30404 = n12128 & n30403;
  assign n30405 = n12157 & n30404;
  assign n30406 = ~n30393 & ~n30405;
  assign n30407 = pi204 & ~n10939;
  assign n30408 = n12473 & n30407;
  assign n30409 = n12317 & n30408;
  assign n30410 = n12316 & n30409;
  assign n30411 = ~n11188 & n30410;
  assign n30412 = ~n12314 & n30411;
  assign n30413 = ~n11510 & n30412;
  assign n30414 = ~n11505 & n30413;
  assign n30415 = n11970 & n30414;
  assign n30416 = n12325 & n30415;
  assign n30417 = n12313 & n30416;
  assign n30418 = n12379 & n30417;
  assign n30419 = n5062 & n28036;
  assign n30420 = n11861 & n30419;
  assign n30421 = ~n3940 & n30420;
  assign n30422 = ~n4001 & n30421;
  assign n30423 = ~n5043 & n30422;
  assign n30424 = ~n5943 & n30423;
  assign n30425 = ~n6951 & n30424;
  assign n30426 = ~n8037 & n30425;
  assign n30427 = ~n9200 & n30426;
  assign n30428 = ~n11813 & n30427;
  assign n30429 = ~n11812 & n30428;
  assign n30430 = ~n11510 & n30429;
  assign n30431 = ~n10445 & n30430;
  assign n30432 = ~n11811 & n30431;
  assign n30433 = n11810 & n30432;
  assign n30434 = n11805 & n30433;
  assign n30435 = n11845 & n30434;
  assign n30436 = ~n30418 & ~n30435;
  assign n30437 = n30406 & n30436;
  assign n30438 = ~n9533 & n27859;
  assign n30439 = ~n11510 & n30438;
  assign n30440 = ~n10787 & n30439;
  assign n30441 = ~n11478 & n30440;
  assign n30442 = n11593 & n30441;
  assign n30443 = n11508 & n30442;
  assign n30444 = n11610 & n30443;
  assign n30445 = n7177 & n28055;
  assign n30446 = n8261 & n30445;
  assign n30447 = ~n6784 & n30446;
  assign n30448 = ~n7158 & n30447;
  assign n30449 = ~n8250 & n30448;
  assign n30450 = ~n9414 & n30449;
  assign n30451 = ~n12053 & n30450;
  assign n30452 = ~n12052 & n30451;
  assign n30453 = ~n11510 & n30452;
  assign n30454 = ~n10667 & n30453;
  assign n30455 = ~n12051 & n30454;
  assign n30456 = n11508 & n30455;
  assign n30457 = n12050 & n30456;
  assign n30458 = n12082 & n30457;
  assign n30459 = ~n30444 & ~n30458;
  assign n30460 = ~n10094 & n27867;
  assign n30461 = ~n11510 & n30460;
  assign n30462 = ~n11318 & n30461;
  assign n30463 = ~n11501 & n30462;
  assign n30464 = n11508 & n30463;
  assign n30465 = n12175 & n30464;
  assign n30466 = n12168 & n30465;
  assign n30467 = ~n9453 & n27990;
  assign n30468 = ~n11510 & n30467;
  assign n30469 = ~n10705 & n30468;
  assign n30470 = ~n12112 & n30469;
  assign n30471 = n12118 & n30470;
  assign n30472 = n11508 & n30471;
  assign n30473 = n12111 & n30472;
  assign n30474 = ~n30466 & ~n30473;
  assign n30475 = n30459 & n30474;
  assign n30476 = n30437 & n30475;
  assign n30477 = n30385 & n30476;
  assign po117 = ~n30329 | ~n30477;
  assign n30479 = ~n10460 & n28153;
  assign n30480 = ~n11510 & n30479;
  assign n30481 = ~n11852 & n30480;
  assign n30482 = n11859 & n30481;
  assign n30483 = ~n10400 & n28157;
  assign n30484 = ~n11790 & n30483;
  assign n30485 = n11795 & n30484;
  assign n30486 = pi229 & ~n501;
  assign n30487 = n12872 & n30486;
  assign n30488 = n14253 & n30487;
  assign n30489 = n12564 & n30488;
  assign n30490 = n28654 & n30489;
  assign n30491 = n12548 & n30490;
  assign n30492 = ~n1172 & n30491;
  assign n30493 = ~n996 & n30492;
  assign n30494 = ~n2306 & n30493;
  assign n30495 = n12571 & n30494;
  assign n30496 = n6677 & n30495;
  assign n30497 = n12580 & n30496;
  assign n30498 = n28668 & n30497;
  assign n30499 = n12542 & n30498;
  assign n30500 = n28650 & n30499;
  assign n30501 = ~n7236 & n30500;
  assign n30502 = ~n6137 & n30501;
  assign n30503 = n6193 & n30502;
  assign n30504 = n6134 & n30503;
  assign n30505 = ~n8867 & n30504;
  assign n30506 = ~n7235 & n30505;
  assign n30507 = n7296 & n30506;
  assign n30508 = n7231 & n30507;
  assign n30509 = ~n10027 & n30508;
  assign n30510 = ~n8866 & n30509;
  assign n30511 = n8898 & n30510;
  assign n30512 = n8863 & n30511;
  assign n30513 = pi221 & ~n501;
  assign n30514 = n12611 & n30513;
  assign n30515 = n26571 & n30514;
  assign n30516 = n12619 & n30515;
  assign n30517 = n28689 & n30516;
  assign n30518 = n12601 & n30517;
  assign n30519 = ~n1172 & n30518;
  assign n30520 = ~n996 & n30519;
  assign n30521 = ~n2306 & n30520;
  assign n30522 = n12626 & n30521;
  assign n30523 = n12628 & n30522;
  assign n30524 = n3823 & n30523;
  assign n30525 = n12634 & n30524;
  assign n30526 = n12682 & n30525;
  assign n30527 = n12844 & n30526;
  assign n30528 = ~n7236 & n30527;
  assign n30529 = ~n6137 & n30528;
  assign n30530 = n6193 & n30529;
  assign n30531 = n6134 & n30530;
  assign n30532 = ~n8867 & n30531;
  assign n30533 = ~n7235 & n30532;
  assign n30534 = n7296 & n30533;
  assign n30535 = n7231 & n30534;
  assign n30536 = ~n10027 & n30535;
  assign n30537 = ~n8866 & n30536;
  assign n30538 = n8898 & n30537;
  assign n30539 = n8863 & n30538;
  assign n30540 = ~n30512 & ~n30539;
  assign n30541 = ~n10788 & ~n30540;
  assign n30542 = ~n10026 & n30541;
  assign n30543 = n10072 & n30542;
  assign n30544 = n10021 & n30543;
  assign n30545 = ~n30485 & ~n30544;
  assign n30546 = ~n30482 & n30545;
  assign n30547 = ~n10554 & n28219;
  assign n30548 = ~n11510 & n30547;
  assign n30549 = ~n11506 & n30548;
  assign n30550 = n11957 & n30549;
  assign n30551 = n11952 & n30550;
  assign n30552 = ~n10629 & n28224;
  assign n30553 = ~n11510 & n30552;
  assign n30554 = n11970 & n30553;
  assign n30555 = n12039 & n30554;
  assign n30556 = n12034 & n30555;
  assign n30557 = ~n30551 & ~n30556;
  assign n30558 = n30546 & n30557;
  assign n30559 = n12275 & n28140;
  assign n30560 = n11562 & n30559;
  assign n30561 = n11560 & n30560;
  assign n30562 = ~n9929 & n30561;
  assign n30563 = ~n11558 & n30562;
  assign n30564 = ~n11557 & n30563;
  assign n30565 = ~n11510 & n30564;
  assign n30566 = ~n11266 & n30565;
  assign n30567 = ~n11509 & n30566;
  assign n30568 = n11508 & n30567;
  assign n30569 = n11556 & n30568;
  assign n30570 = n11587 & n30569;
  assign n30571 = n11681 & n28263;
  assign n30572 = n11680 & n30571;
  assign n30573 = ~n1372 & n30572;
  assign n30574 = ~n2243 & n30573;
  assign n30575 = ~n3104 & n30574;
  assign n30576 = ~n3971 & n30575;
  assign n30577 = ~n4003 & n30576;
  assign n30578 = ~n4872 & n30577;
  assign n30579 = ~n5801 & n30578;
  assign n30580 = ~n6739 & n30579;
  assign n30581 = ~n7807 & n30580;
  assign n30582 = ~n8989 & n30581;
  assign n30583 = ~n10273 & n30582;
  assign n30584 = ~n11678 & n30583;
  assign n30585 = ~n11677 & n30584;
  assign n30586 = ~n11676 & n30585;
  assign n30587 = ~n11499 & n30586;
  assign n30588 = ~n11675 & n30587;
  assign n30589 = n11674 & n30588;
  assign n30590 = n11669 & n30589;
  assign n30591 = n11716 & n30590;
  assign n30592 = ~n30570 & ~n30591;
  assign n30593 = pi061 & ~n2176;
  assign n30594 = n4955 & n30593;
  assign n30595 = n7909 & n30594;
  assign n30596 = ~n2242 & n30595;
  assign n30597 = ~n3095 & n30596;
  assign n30598 = ~n3997 & n30597;
  assign n30599 = ~n4003 & n30598;
  assign n30600 = ~n4837 & n30599;
  assign n30601 = ~n5822 & n30600;
  assign n30602 = ~n6820 & n30601;
  assign n30603 = ~n7785 & n30602;
  assign n30604 = ~n9027 & n30603;
  assign n30605 = ~n10245 & n30604;
  assign n30606 = ~n11733 & n30605;
  assign n30607 = ~n11732 & n30606;
  assign n30608 = ~n11731 & n30607;
  assign n30609 = ~n11536 & n30608;
  assign n30610 = ~n11730 & n30609;
  assign n30611 = n11729 & n30610;
  assign n30612 = n11724 & n30611;
  assign n30613 = n11768 & n30612;
  assign n30614 = n12013 & n22732;
  assign n30615 = ~n5808 & n30614;
  assign n30616 = ~n6056 & n30615;
  assign n30617 = ~n7073 & n30616;
  assign n30618 = ~n8179 & n30617;
  assign n30619 = ~n9344 & n30618;
  assign n30620 = ~n11974 & n30619;
  assign n30621 = ~n11973 & n30620;
  assign n30622 = ~n11510 & n30621;
  assign n30623 = ~n10594 & n30622;
  assign n30624 = ~n11972 & n30623;
  assign n30625 = n11971 & n30624;
  assign n30626 = n11968 & n30625;
  assign n30627 = n12004 & n30626;
  assign n30628 = ~n30613 & ~n30627;
  assign n30629 = n30592 & n30628;
  assign n30630 = n30558 & n30629;
  assign n30631 = n5085 & n28335;
  assign n30632 = n11931 & n30631;
  assign n30633 = ~n4817 & n30632;
  assign n30634 = ~n4902 & n30633;
  assign n30635 = ~n6001 & n30634;
  assign n30636 = ~n7014 & n30635;
  assign n30637 = ~n8114 & n30636;
  assign n30638 = ~n9276 & n30637;
  assign n30639 = ~n11898 & n30638;
  assign n30640 = ~n11897 & n30639;
  assign n30641 = ~n11510 & n30640;
  assign n30642 = ~n10523 & n30641;
  assign n30643 = ~n11896 & n30642;
  assign n30644 = n11895 & n30643;
  assign n30645 = n11891 & n30644;
  assign n30646 = n11927 & n30645;
  assign n30647 = n11378 & n26066;
  assign n30648 = n9942 & n30647;
  assign n30649 = ~n8834 & n30648;
  assign n30650 = ~n10002 & n30649;
  assign n30651 = ~n12212 & n30650;
  assign n30652 = ~n12211 & n30651;
  assign n30653 = ~n11510 & n30652;
  assign n30654 = ~n11297 & n30653;
  assign n30655 = ~n11478 & n30654;
  assign n30656 = n11508 & n30655;
  assign n30657 = n12210 & n30656;
  assign n30658 = n12239 & n30657;
  assign n30659 = ~n30646 & ~n30658;
  assign n30660 = n9115 & n22782;
  assign n30661 = ~n3066 & n30660;
  assign n30662 = ~n3983 & n30661;
  assign n30663 = ~n4003 & n30662;
  assign n30664 = ~n4024 & n30663;
  assign n30665 = ~n4999 & n30664;
  assign n30666 = ~n5827 & n30665;
  assign n30667 = ~n6893 & n30666;
  assign n30668 = ~n7890 & n30667;
  assign n30669 = ~n9131 & n30668;
  assign n30670 = ~n11627 & n30669;
  assign n30671 = ~n11626 & n30670;
  assign n30672 = ~n11625 & n30671;
  assign n30673 = ~n10278 & n30672;
  assign n30674 = ~n11624 & n30673;
  assign n30675 = n11623 & n30674;
  assign n30676 = n11618 & n30675;
  assign n30677 = n11661 & n30676;
  assign n30678 = pi197 & ~n10074;
  assign n30679 = ~n11510 & n30678;
  assign n30680 = ~n11343 & n30679;
  assign n30681 = ~n11509 & n30680;
  assign n30682 = n11508 & n30681;
  assign n30683 = n11503 & n30682;
  assign n30684 = n11550 & n30683;
  assign n30685 = ~n30677 & ~n30684;
  assign n30686 = n30659 & n30685;
  assign n30687 = pi213 & ~n10879;
  assign n30688 = ~n12412 & n30687;
  assign n30689 = ~n11510 & n30688;
  assign n30690 = ~n11505 & n30689;
  assign n30691 = n11970 & n30690;
  assign n30692 = n12325 & n30691;
  assign n30693 = n12411 & n30692;
  assign n30694 = n12470 & n30693;
  assign n30695 = n12182 & n24400;
  assign n30696 = ~n7869 & n30695;
  assign n30697 = ~n8346 & n30696;
  assign n30698 = ~n9485 & n30697;
  assign n30699 = ~n12130 & n30698;
  assign n30700 = ~n12129 & n30699;
  assign n30701 = ~n11510 & n30700;
  assign n30702 = ~n10741 & n30701;
  assign n30703 = ~n11501 & n30702;
  assign n30704 = n11508 & n30703;
  assign n30705 = n12128 & n30704;
  assign n30706 = n12157 & n30705;
  assign n30707 = ~n30694 & ~n30706;
  assign n30708 = pi205 & ~n10939;
  assign n30709 = n12473 & n30708;
  assign n30710 = n12317 & n30709;
  assign n30711 = n12316 & n30710;
  assign n30712 = ~n11188 & n30711;
  assign n30713 = ~n12314 & n30712;
  assign n30714 = ~n11510 & n30713;
  assign n30715 = ~n11505 & n30714;
  assign n30716 = n11970 & n30715;
  assign n30717 = n12325 & n30716;
  assign n30718 = n12313 & n30717;
  assign n30719 = n12379 & n30718;
  assign n30720 = n5062 & n28302;
  assign n30721 = n11861 & n30720;
  assign n30722 = ~n3940 & n30721;
  assign n30723 = ~n4001 & n30722;
  assign n30724 = ~n5043 & n30723;
  assign n30725 = ~n5943 & n30724;
  assign n30726 = ~n6951 & n30725;
  assign n30727 = ~n8037 & n30726;
  assign n30728 = ~n9200 & n30727;
  assign n30729 = ~n11813 & n30728;
  assign n30730 = ~n11812 & n30729;
  assign n30731 = ~n11510 & n30730;
  assign n30732 = ~n10445 & n30731;
  assign n30733 = ~n11811 & n30732;
  assign n30734 = n11810 & n30733;
  assign n30735 = n11805 & n30734;
  assign n30736 = n11845 & n30735;
  assign n30737 = ~n30719 & ~n30736;
  assign n30738 = n30707 & n30737;
  assign n30739 = ~n9533 & n28125;
  assign n30740 = ~n11510 & n30739;
  assign n30741 = ~n10787 & n30740;
  assign n30742 = ~n11478 & n30741;
  assign n30743 = n11593 & n30742;
  assign n30744 = n11508 & n30743;
  assign n30745 = n11610 & n30744;
  assign n30746 = n7177 & n28321;
  assign n30747 = n8261 & n30746;
  assign n30748 = ~n6784 & n30747;
  assign n30749 = ~n7158 & n30748;
  assign n30750 = ~n8250 & n30749;
  assign n30751 = ~n9414 & n30750;
  assign n30752 = ~n12053 & n30751;
  assign n30753 = ~n12052 & n30752;
  assign n30754 = ~n11510 & n30753;
  assign n30755 = ~n10667 & n30754;
  assign n30756 = ~n12051 & n30755;
  assign n30757 = n11508 & n30756;
  assign n30758 = n12050 & n30757;
  assign n30759 = n12082 & n30758;
  assign n30760 = ~n30745 & ~n30759;
  assign n30761 = ~n10094 & n28133;
  assign n30762 = ~n11510 & n30761;
  assign n30763 = ~n11318 & n30762;
  assign n30764 = ~n11501 & n30763;
  assign n30765 = n11508 & n30764;
  assign n30766 = n12175 & n30765;
  assign n30767 = n12168 & n30766;
  assign n30768 = ~n9453 & n28256;
  assign n30769 = ~n11510 & n30768;
  assign n30770 = ~n10705 & n30769;
  assign n30771 = ~n12112 & n30770;
  assign n30772 = n12118 & n30771;
  assign n30773 = n11508 & n30772;
  assign n30774 = n12111 & n30773;
  assign n30775 = ~n30767 & ~n30774;
  assign n30776 = n30760 & n30775;
  assign n30777 = n30738 & n30776;
  assign n30778 = n30686 & n30777;
  assign po118 = ~n30630 | ~n30778;
  assign n30780 = ~n10460 & n28419;
  assign n30781 = ~n11510 & n30780;
  assign n30782 = ~n11852 & n30781;
  assign n30783 = n11859 & n30782;
  assign n30784 = ~n10400 & n28423;
  assign n30785 = ~n11790 & n30784;
  assign n30786 = n11795 & n30785;
  assign n30787 = pi230 & ~n501;
  assign n30788 = n12872 & n30787;
  assign n30789 = n14253 & n30788;
  assign n30790 = n12564 & n30789;
  assign n30791 = n28654 & n30790;
  assign n30792 = n12548 & n30791;
  assign n30793 = ~n1172 & n30792;
  assign n30794 = ~n996 & n30793;
  assign n30795 = ~n2306 & n30794;
  assign n30796 = n12571 & n30795;
  assign n30797 = n6677 & n30796;
  assign n30798 = n12580 & n30797;
  assign n30799 = n28668 & n30798;
  assign n30800 = n12542 & n30799;
  assign n30801 = n28650 & n30800;
  assign n30802 = ~n7236 & n30801;
  assign n30803 = ~n6137 & n30802;
  assign n30804 = n6193 & n30803;
  assign n30805 = n6134 & n30804;
  assign n30806 = ~n8867 & n30805;
  assign n30807 = ~n7235 & n30806;
  assign n30808 = n7296 & n30807;
  assign n30809 = n7231 & n30808;
  assign n30810 = ~n10027 & n30809;
  assign n30811 = ~n8866 & n30810;
  assign n30812 = n8898 & n30811;
  assign n30813 = n8863 & n30812;
  assign n30814 = pi222 & ~n501;
  assign n30815 = n12611 & n30814;
  assign n30816 = n26571 & n30815;
  assign n30817 = n12619 & n30816;
  assign n30818 = n28689 & n30817;
  assign n30819 = n12601 & n30818;
  assign n30820 = ~n1172 & n30819;
  assign n30821 = ~n996 & n30820;
  assign n30822 = ~n2306 & n30821;
  assign n30823 = n12626 & n30822;
  assign n30824 = n12628 & n30823;
  assign n30825 = n3823 & n30824;
  assign n30826 = n12634 & n30825;
  assign n30827 = n12682 & n30826;
  assign n30828 = n12844 & n30827;
  assign n30829 = ~n7236 & n30828;
  assign n30830 = ~n6137 & n30829;
  assign n30831 = n6193 & n30830;
  assign n30832 = n6134 & n30831;
  assign n30833 = ~n8867 & n30832;
  assign n30834 = ~n7235 & n30833;
  assign n30835 = n7296 & n30834;
  assign n30836 = n7231 & n30835;
  assign n30837 = ~n10027 & n30836;
  assign n30838 = ~n8866 & n30837;
  assign n30839 = n8898 & n30838;
  assign n30840 = n8863 & n30839;
  assign n30841 = ~n30813 & ~n30840;
  assign n30842 = ~n10788 & ~n30841;
  assign n30843 = ~n10026 & n30842;
  assign n30844 = n10072 & n30843;
  assign n30845 = n10021 & n30844;
  assign n30846 = ~n30786 & ~n30845;
  assign n30847 = ~n30783 & n30846;
  assign n30848 = ~n10554 & n28485;
  assign n30849 = ~n11510 & n30848;
  assign n30850 = ~n11506 & n30849;
  assign n30851 = n11957 & n30850;
  assign n30852 = n11952 & n30851;
  assign n30853 = ~n10629 & n28490;
  assign n30854 = ~n11510 & n30853;
  assign n30855 = n11970 & n30854;
  assign n30856 = n12039 & n30855;
  assign n30857 = n12034 & n30856;
  assign n30858 = ~n30852 & ~n30857;
  assign n30859 = n30847 & n30858;
  assign n30860 = n12275 & n28406;
  assign n30861 = n11562 & n30860;
  assign n30862 = n11560 & n30861;
  assign n30863 = ~n9929 & n30862;
  assign n30864 = ~n11558 & n30863;
  assign n30865 = ~n11557 & n30864;
  assign n30866 = ~n11510 & n30865;
  assign n30867 = ~n11266 & n30866;
  assign n30868 = ~n11509 & n30867;
  assign n30869 = n11508 & n30868;
  assign n30870 = n11556 & n30869;
  assign n30871 = n11587 & n30870;
  assign n30872 = n11681 & n28529;
  assign n30873 = n11680 & n30872;
  assign n30874 = ~n1372 & n30873;
  assign n30875 = ~n2243 & n30874;
  assign n30876 = ~n3104 & n30875;
  assign n30877 = ~n3971 & n30876;
  assign n30878 = ~n4003 & n30877;
  assign n30879 = ~n4872 & n30878;
  assign n30880 = ~n5801 & n30879;
  assign n30881 = ~n6739 & n30880;
  assign n30882 = ~n7807 & n30881;
  assign n30883 = ~n8989 & n30882;
  assign n30884 = ~n10273 & n30883;
  assign n30885 = ~n11678 & n30884;
  assign n30886 = ~n11677 & n30885;
  assign n30887 = ~n11676 & n30886;
  assign n30888 = ~n11499 & n30887;
  assign n30889 = ~n11675 & n30888;
  assign n30890 = n11674 & n30889;
  assign n30891 = n11669 & n30890;
  assign n30892 = n11716 & n30891;
  assign n30893 = ~n30871 & ~n30892;
  assign n30894 = pi062 & ~n2176;
  assign n30895 = n4955 & n30894;
  assign n30896 = n7909 & n30895;
  assign n30897 = ~n2242 & n30896;
  assign n30898 = ~n3095 & n30897;
  assign n30899 = ~n3997 & n30898;
  assign n30900 = ~n4003 & n30899;
  assign n30901 = ~n4837 & n30900;
  assign n30902 = ~n5822 & n30901;
  assign n30903 = ~n6820 & n30902;
  assign n30904 = ~n7785 & n30903;
  assign n30905 = ~n9027 & n30904;
  assign n30906 = ~n10245 & n30905;
  assign n30907 = ~n11733 & n30906;
  assign n30908 = ~n11732 & n30907;
  assign n30909 = ~n11731 & n30908;
  assign n30910 = ~n11536 & n30909;
  assign n30911 = ~n11730 & n30910;
  assign n30912 = n11729 & n30911;
  assign n30913 = n11724 & n30912;
  assign n30914 = n11768 & n30913;
  assign n30915 = n12013 & n22899;
  assign n30916 = ~n5808 & n30915;
  assign n30917 = ~n6056 & n30916;
  assign n30918 = ~n7073 & n30917;
  assign n30919 = ~n8179 & n30918;
  assign n30920 = ~n9344 & n30919;
  assign n30921 = ~n11974 & n30920;
  assign n30922 = ~n11973 & n30921;
  assign n30923 = ~n11510 & n30922;
  assign n30924 = ~n10594 & n30923;
  assign n30925 = ~n11972 & n30924;
  assign n30926 = n11971 & n30925;
  assign n30927 = n11968 & n30926;
  assign n30928 = n12004 & n30927;
  assign n30929 = ~n30914 & ~n30928;
  assign n30930 = n30893 & n30929;
  assign n30931 = n30859 & n30930;
  assign n30932 = n5085 & n28601;
  assign n30933 = n11931 & n30932;
  assign n30934 = ~n4817 & n30933;
  assign n30935 = ~n4902 & n30934;
  assign n30936 = ~n6001 & n30935;
  assign n30937 = ~n7014 & n30936;
  assign n30938 = ~n8114 & n30937;
  assign n30939 = ~n9276 & n30938;
  assign n30940 = ~n11898 & n30939;
  assign n30941 = ~n11897 & n30940;
  assign n30942 = ~n11510 & n30941;
  assign n30943 = ~n10523 & n30942;
  assign n30944 = ~n11896 & n30943;
  assign n30945 = n11895 & n30944;
  assign n30946 = n11891 & n30945;
  assign n30947 = n11927 & n30946;
  assign n30948 = n11378 & n26299;
  assign n30949 = n9942 & n30948;
  assign n30950 = ~n8834 & n30949;
  assign n30951 = ~n10002 & n30950;
  assign n30952 = ~n12212 & n30951;
  assign n30953 = ~n12211 & n30952;
  assign n30954 = ~n11510 & n30953;
  assign n30955 = ~n11297 & n30954;
  assign n30956 = ~n11478 & n30955;
  assign n30957 = n11508 & n30956;
  assign n30958 = n12210 & n30957;
  assign n30959 = n12239 & n30958;
  assign n30960 = ~n30947 & ~n30959;
  assign n30961 = n9115 & n22949;
  assign n30962 = ~n3066 & n30961;
  assign n30963 = ~n3983 & n30962;
  assign n30964 = ~n4003 & n30963;
  assign n30965 = ~n4024 & n30964;
  assign n30966 = ~n4999 & n30965;
  assign n30967 = ~n5827 & n30966;
  assign n30968 = ~n6893 & n30967;
  assign n30969 = ~n7890 & n30968;
  assign n30970 = ~n9131 & n30969;
  assign n30971 = ~n11627 & n30970;
  assign n30972 = ~n11626 & n30971;
  assign n30973 = ~n11625 & n30972;
  assign n30974 = ~n10278 & n30973;
  assign n30975 = ~n11624 & n30974;
  assign n30976 = n11623 & n30975;
  assign n30977 = n11618 & n30976;
  assign n30978 = n11661 & n30977;
  assign n30979 = pi198 & ~n10074;
  assign n30980 = ~n11510 & n30979;
  assign n30981 = ~n11343 & n30980;
  assign n30982 = ~n11509 & n30981;
  assign n30983 = n11508 & n30982;
  assign n30984 = n11503 & n30983;
  assign n30985 = n11550 & n30984;
  assign n30986 = ~n30978 & ~n30985;
  assign n30987 = n30960 & n30986;
  assign n30988 = pi214 & ~n10879;
  assign n30989 = ~n12412 & n30988;
  assign n30990 = ~n11510 & n30989;
  assign n30991 = ~n11505 & n30990;
  assign n30992 = n11970 & n30991;
  assign n30993 = n12325 & n30992;
  assign n30994 = n12411 & n30993;
  assign n30995 = n12470 & n30994;
  assign n30996 = n12182 & n24593;
  assign n30997 = ~n7869 & n30996;
  assign n30998 = ~n8346 & n30997;
  assign n30999 = ~n9485 & n30998;
  assign n31000 = ~n12130 & n30999;
  assign n31001 = ~n12129 & n31000;
  assign n31002 = ~n11510 & n31001;
  assign n31003 = ~n10741 & n31002;
  assign n31004 = ~n11501 & n31003;
  assign n31005 = n11508 & n31004;
  assign n31006 = n12128 & n31005;
  assign n31007 = n12157 & n31006;
  assign n31008 = ~n30995 & ~n31007;
  assign n31009 = pi206 & ~n10939;
  assign n31010 = n12473 & n31009;
  assign n31011 = n12317 & n31010;
  assign n31012 = n12316 & n31011;
  assign n31013 = ~n11188 & n31012;
  assign n31014 = ~n12314 & n31013;
  assign n31015 = ~n11510 & n31014;
  assign n31016 = ~n11505 & n31015;
  assign n31017 = n11970 & n31016;
  assign n31018 = n12325 & n31017;
  assign n31019 = n12313 & n31018;
  assign n31020 = n12379 & n31019;
  assign n31021 = n5062 & n28568;
  assign n31022 = n11861 & n31021;
  assign n31023 = ~n3940 & n31022;
  assign n31024 = ~n4001 & n31023;
  assign n31025 = ~n5043 & n31024;
  assign n31026 = ~n5943 & n31025;
  assign n31027 = ~n6951 & n31026;
  assign n31028 = ~n8037 & n31027;
  assign n31029 = ~n9200 & n31028;
  assign n31030 = ~n11813 & n31029;
  assign n31031 = ~n11812 & n31030;
  assign n31032 = ~n11510 & n31031;
  assign n31033 = ~n10445 & n31032;
  assign n31034 = ~n11811 & n31033;
  assign n31035 = n11810 & n31034;
  assign n31036 = n11805 & n31035;
  assign n31037 = n11845 & n31036;
  assign n31038 = ~n31020 & ~n31037;
  assign n31039 = n31008 & n31038;
  assign n31040 = ~n9533 & n28391;
  assign n31041 = ~n11510 & n31040;
  assign n31042 = ~n10787 & n31041;
  assign n31043 = ~n11478 & n31042;
  assign n31044 = n11593 & n31043;
  assign n31045 = n11508 & n31044;
  assign n31046 = n11610 & n31045;
  assign n31047 = n7177 & n28587;
  assign n31048 = n8261 & n31047;
  assign n31049 = ~n6784 & n31048;
  assign n31050 = ~n7158 & n31049;
  assign n31051 = ~n8250 & n31050;
  assign n31052 = ~n9414 & n31051;
  assign n31053 = ~n12053 & n31052;
  assign n31054 = ~n12052 & n31053;
  assign n31055 = ~n11510 & n31054;
  assign n31056 = ~n10667 & n31055;
  assign n31057 = ~n12051 & n31056;
  assign n31058 = n11508 & n31057;
  assign n31059 = n12050 & n31058;
  assign n31060 = n12082 & n31059;
  assign n31061 = ~n31046 & ~n31060;
  assign n31062 = ~n10094 & n28399;
  assign n31063 = ~n11510 & n31062;
  assign n31064 = ~n11318 & n31063;
  assign n31065 = ~n11501 & n31064;
  assign n31066 = n11508 & n31065;
  assign n31067 = n12175 & n31066;
  assign n31068 = n12168 & n31067;
  assign n31069 = ~n9453 & n28522;
  assign n31070 = ~n11510 & n31069;
  assign n31071 = ~n10705 & n31070;
  assign n31072 = ~n12112 & n31071;
  assign n31073 = n12118 & n31072;
  assign n31074 = n11508 & n31073;
  assign n31075 = n12111 & n31074;
  assign n31076 = ~n31068 & ~n31075;
  assign n31077 = n31061 & n31076;
  assign n31078 = n31039 & n31077;
  assign n31079 = n30987 & n31078;
  assign po119 = ~n30931 | ~n31079;
  assign n31081 = ~n10705 & n28792;
  assign n31082 = ~n12861 & n31081;
  assign n31083 = ~n12121 & n31082;
  assign n31084 = ~n13717 & n31083;
  assign n31085 = n13723 & n31084;
  assign n31086 = n13095 & n31085;
  assign n31087 = n13716 & n31086;
  assign n31088 = ~n11318 & n28841;
  assign n31089 = ~n12861 & n31088;
  assign n31090 = ~n12181 & n31089;
  assign n31091 = ~n13052 & n31090;
  assign n31092 = n13095 & n31091;
  assign n31093 = n13758 & n31092;
  assign n31094 = n13751 & n31093;
  assign n31095 = ~n31087 & ~n31094;
  assign n31096 = ~n10787 & n28808;
  assign n31097 = ~n12861 & n31096;
  assign n31098 = ~n11611 & n31097;
  assign n31099 = ~n12973 & n31098;
  assign n31100 = n13802 & n31099;
  assign n31101 = n13095 & n31100;
  assign n31102 = n13819 & n31101;
  assign n31103 = ~n11343 & n28768;
  assign n31104 = ~n12861 & n31103;
  assign n31105 = ~n11551 & n31104;
  assign n31106 = ~n12973 & n31105;
  assign n31107 = n13095 & n31106;
  assign n31108 = n13885 & n31107;
  assign n31109 = n13905 & n31108;
  assign n31110 = ~n31102 & ~n31109;
  assign n31111 = n31095 & n31110;
  assign n31112 = pi039 & ~n1204;
  assign n31113 = ~n776 & ~n1205;
  assign n31114 = ~n777 & n31113;
  assign n31115 = n31112 & n31114;
  assign n31116 = ~n1203 & n31115;
  assign n31117 = ~n775 & n31116;
  assign n31118 = ~n1238 & n31117;
  assign n31119 = ~n688 & ~n750;
  assign n31120 = ~n718 & n31119;
  assign n31121 = n31118 & n31120;
  assign n31122 = ~n1372 & n31121;
  assign n31123 = ~n2243 & n31122;
  assign n31124 = ~n3104 & n31123;
  assign n31125 = ~n3971 & n31124;
  assign n31126 = ~n4003 & n31125;
  assign n31127 = ~n4872 & n31126;
  assign n31128 = ~n5801 & n31127;
  assign n31129 = ~n6739 & n31128;
  assign n31130 = ~n7807 & n31129;
  assign n31131 = ~n8989 & n31130;
  assign n31132 = ~n10273 & n31131;
  assign n31133 = ~n13200 & n31132;
  assign n31134 = ~n13199 & n31133;
  assign n31135 = ~n11499 & n31134;
  assign n31136 = ~n13198 & n31135;
  assign n31137 = ~n13076 & n31136;
  assign n31138 = ~n13197 & n31137;
  assign n31139 = n13223 & n31138;
  assign n31140 = n13196 & n31139;
  assign n31141 = n13248 & n31140;
  assign n31142 = ~n11860 & n28729;
  assign n31143 = ~n12861 & n31142;
  assign n31144 = ~n13399 & n31143;
  assign n31145 = n13406 & n31144;
  assign n31146 = ~n13312 & n28644;
  assign n31147 = ~n13310 & n31146;
  assign n31148 = n13317 & n31147;
  assign n31149 = pi231 & ~n501;
  assign n31150 = n14255 & n31149;
  assign n31151 = n14253 & n31150;
  assign n31152 = n14261 & n14487;
  assign n31153 = n5716 & n31152;
  assign n31154 = n14260 & n31153;
  assign n31155 = n31151 & n31154;
  assign n31156 = ~n3285 & ~n3375;
  assign n31157 = n4796 & n31156;
  assign n31158 = n14275 & n31157;
  assign n31159 = n5720 & n12550;
  assign n31160 = n14278 & n31159;
  assign n31161 = n31158 & n31160;
  assign n31162 = n14274 & n31161;
  assign n31163 = n31155 & n31162;
  assign n31164 = ~n1172 & n31163;
  assign n31165 = ~n996 & n31164;
  assign n31166 = ~n2306 & n31165;
  assign n31167 = n3819 & n31166;
  assign n31168 = n14139 & n31167;
  assign n31169 = n12583 & n31168;
  assign n31170 = n14252 & n31169;
  assign n31171 = n14242 & n31170;
  assign n31172 = n14431 & n31171;
  assign n31173 = ~n7236 & n31172;
  assign n31174 = ~n6137 & n31173;
  assign n31175 = n6193 & n31174;
  assign n31176 = n6134 & n31175;
  assign n31177 = ~n8867 & n31176;
  assign n31178 = ~n7235 & n31177;
  assign n31179 = n7296 & n31178;
  assign n31180 = n7231 & n31179;
  assign n31181 = ~n10027 & n31180;
  assign n31182 = ~n8866 & n31181;
  assign n31183 = n8898 & n31182;
  assign n31184 = n8863 & n31183;
  assign n31185 = pi239 & ~n501;
  assign n31186 = n14188 & n31185;
  assign n31187 = n14194 & n14536;
  assign n31188 = n14197 & n31187;
  assign n31189 = n14193 & n31188;
  assign n31190 = n31186 & n31189;
  assign n31191 = n14210 & n31156;
  assign n31192 = n6142 & n31191;
  assign n31193 = n4796 & n12550;
  assign n31194 = n14539 & n31193;
  assign n31195 = n31192 & n31194;
  assign n31196 = n14209 & n31195;
  assign n31197 = n31190 & n31196;
  assign n31198 = ~n1172 & n31197;
  assign n31199 = ~n996 & n31198;
  assign n31200 = ~n2306 & n31199;
  assign n31201 = n3819 & n31200;
  assign n31202 = n3821 & n31201;
  assign n31203 = n14186 & n31202;
  assign n31204 = n14229 & n31203;
  assign n31205 = n14184 & n31204;
  assign n31206 = n14180 & n31205;
  assign n31207 = ~n7236 & n31206;
  assign n31208 = ~n6137 & n31207;
  assign n31209 = n6193 & n31208;
  assign n31210 = n6134 & n31209;
  assign n31211 = ~n8867 & n31210;
  assign n31212 = ~n7235 & n31211;
  assign n31213 = n7296 & n31212;
  assign n31214 = n7231 & n31213;
  assign n31215 = ~n10027 & n31214;
  assign n31216 = ~n8866 & n31215;
  assign n31217 = n8898 & n31216;
  assign n31218 = n8863 & n31217;
  assign n31219 = ~n31184 & ~n31218;
  assign n31220 = ~n10788 & ~n31219;
  assign n31221 = ~n10026 & n31220;
  assign n31222 = n10072 & n31221;
  assign n31223 = n10021 & n31222;
  assign n31224 = ~n31148 & ~n31223;
  assign n31225 = ~n31145 & n31224;
  assign n31226 = ~n11959 & n28639;
  assign n31227 = ~n12861 & n31226;
  assign n31228 = ~n12950 & n31227;
  assign n31229 = n13491 & n31228;
  assign n31230 = n13486 & n31229;
  assign n31231 = ~n12041 & n28724;
  assign n31232 = ~n12861 & n31231;
  assign n31233 = n13094 & n31232;
  assign n31234 = n13577 & n31233;
  assign n31235 = n13572 & n31234;
  assign n31236 = ~n31230 & ~n31235;
  assign n31237 = n31225 & n31236;
  assign n31238 = ~n31141 & n31237;
  assign n31239 = pi215 & pi255;
  assign n31240 = ~n12709 & n31239;
  assign n31241 = ~n12671 & n31240;
  assign n31242 = ~n12811 & n31241;
  assign n31243 = ~n12773 & n13910;
  assign n31244 = n31242 & n31243;
  assign n31245 = ~n12902 & n31244;
  assign n31246 = ~n13908 & n31245;
  assign n31247 = ~n12861 & n31246;
  assign n31248 = ~n12860 & n31247;
  assign n31249 = n12952 & n31248;
  assign n31250 = n13919 & n31249;
  assign n31251 = n14008 & n31250;
  assign n31252 = pi103 & ~n4426;
  assign n31253 = ~n4427 & n31252;
  assign n31254 = ~n4425 & n31253;
  assign n31255 = ~n4707 & n31254;
  assign n31256 = n4490 & n5083;
  assign n31257 = n31255 & n31256;
  assign n31258 = ~n4817 & n31257;
  assign n31259 = ~n4902 & n31258;
  assign n31260 = ~n6001 & n31259;
  assign n31261 = ~n7014 & n31260;
  assign n31262 = ~n8114 & n31261;
  assign n31263 = ~n9276 & n31262;
  assign n31264 = ~n13438 & n31263;
  assign n31265 = ~n13437 & n31264;
  assign n31266 = ~n10523 & n31265;
  assign n31267 = ~n12861 & n31266;
  assign n31268 = ~n11928 & n31267;
  assign n31269 = ~n13436 & n31268;
  assign n31270 = n13453 & n31269;
  assign n31271 = n13435 & n31270;
  assign n31272 = n13478 & n31271;
  assign n31273 = ~n31251 & ~n31272;
  assign n31274 = n31238 & n31273;
  assign n31275 = n31111 & n31274;
  assign n31276 = pi199 & ~n10909;
  assign n31277 = ~n11168 & n31276;
  assign n31278 = n11135 & n31277;
  assign n31279 = ~n11188 & n31278;
  assign n31280 = ~n14011 & n31279;
  assign n31281 = ~n14010 & n31280;
  assign n31282 = ~n12861 & n31281;
  assign n31283 = ~n12380 & n31282;
  assign n31284 = ~n12972 & n31283;
  assign n31285 = n14020 & n31284;
  assign n31286 = n13095 & n31285;
  assign n31287 = n14044 & n31286;
  assign n31288 = n13654 & n23136;
  assign n31289 = ~n7869 & n31288;
  assign n31290 = ~n8346 & n31289;
  assign n31291 = ~n9485 & n31290;
  assign n31292 = ~n13653 & n31291;
  assign n31293 = ~n13652 & n31292;
  assign n31294 = ~n10741 & n31293;
  assign n31295 = ~n12861 & n31294;
  assign n31296 = ~n12158 & n31295;
  assign n31297 = ~n13052 & n31296;
  assign n31298 = n13667 & n31297;
  assign n31299 = n13095 & n31298;
  assign n31300 = n13692 & n31299;
  assign n31301 = ~n12861 & n28799;
  assign n31302 = ~n12471 & n31301;
  assign n31303 = ~n12972 & n31302;
  assign n31304 = n14020 & n31303;
  assign n31305 = n13095 & n31304;
  assign n31306 = n14072 & n31305;
  assign n31307 = ~n31300 & ~n31306;
  assign n31308 = ~n31287 & n31307;
  assign n31309 = pi223 & ~n12946;
  assign n31310 = ~n12903 & n31309;
  assign n31311 = ~n12861 & n31310;
  assign n31312 = ~n12860 & n31311;
  assign n31313 = n12952 & n31312;
  assign n31314 = n12975 & n31313;
  assign n31315 = n13092 & n31314;
  assign n31316 = pi135 & ~n6313;
  assign n31317 = n7175 & n31316;
  assign n31318 = n13694 & n31317;
  assign n31319 = ~n6784 & n31318;
  assign n31320 = ~n7158 & n31319;
  assign n31321 = ~n8250 & n31320;
  assign n31322 = ~n9414 & n31321;
  assign n31323 = ~n13602 & n31322;
  assign n31324 = ~n13601 & n31323;
  assign n31325 = ~n10667 & n31324;
  assign n31326 = ~n12861 & n31325;
  assign n31327 = ~n12083 & n31326;
  assign n31328 = ~n13600 & n31327;
  assign n31329 = n13618 & n31328;
  assign n31330 = n13095 & n31329;
  assign n31331 = n13643 & n31330;
  assign n31332 = ~n31315 & ~n31331;
  assign n31333 = pi055 & ~n1522;
  assign n31334 = ~n1523 & n31333;
  assign n31335 = ~n1521 & n31334;
  assign n31336 = ~n1679 & n31335;
  assign n31337 = n1741 & n3069;
  assign n31338 = n31336 & n31337;
  assign n31339 = ~n2242 & n31338;
  assign n31340 = ~n3095 & n31339;
  assign n31341 = ~n3997 & n31340;
  assign n31342 = ~n4003 & n31341;
  assign n31343 = ~n4837 & n31342;
  assign n31344 = ~n5822 & n31343;
  assign n31345 = ~n6820 & n31344;
  assign n31346 = ~n7785 & n31345;
  assign n31347 = ~n9027 & n31346;
  assign n31348 = ~n10245 & n31347;
  assign n31349 = ~n13258 & n31348;
  assign n31350 = ~n13257 & n31349;
  assign n31351 = ~n11536 & n31350;
  assign n31352 = ~n13256 & n31351;
  assign n31353 = ~n13036 & n31352;
  assign n31354 = ~n13255 & n31353;
  assign n31355 = n13281 & n31354;
  assign n31356 = n13254 & n31355;
  assign n31357 = n13306 & n31356;
  assign n31358 = pi087 & ~n3587;
  assign n31359 = ~n3588 & n31358;
  assign n31360 = ~n3586 & n31359;
  assign n31361 = ~n3710 & n31360;
  assign n31362 = n4096 & n4103;
  assign n31363 = n31361 & n31362;
  assign n31364 = ~n3940 & n31363;
  assign n31365 = ~n4001 & n31364;
  assign n31366 = ~n5043 & n31365;
  assign n31367 = ~n5943 & n31366;
  assign n31368 = ~n6951 & n31367;
  assign n31369 = ~n8037 & n31368;
  assign n31370 = ~n9200 & n31369;
  assign n31371 = ~n13348 & n31370;
  assign n31372 = ~n13347 & n31371;
  assign n31373 = ~n10445 & n31372;
  assign n31374 = ~n12861 & n31373;
  assign n31375 = ~n11846 & n31374;
  assign n31376 = ~n13346 & n31375;
  assign n31377 = n13367 & n31376;
  assign n31378 = n13345 & n31377;
  assign n31379 = n13392 & n31378;
  assign n31380 = ~n31357 & ~n31379;
  assign n31381 = n31332 & n31380;
  assign n31382 = pi167 & ~n8629;
  assign n31383 = ~n8630 & n31382;
  assign n31384 = ~n8628 & n31383;
  assign n31385 = ~n8574 & n31384;
  assign n31386 = n8545 & n31385;
  assign n31387 = ~n8834 & n31386;
  assign n31388 = ~n10002 & n31387;
  assign n31389 = ~n13097 & n31388;
  assign n31390 = ~n13096 & n31389;
  assign n31391 = ~n11297 & n31390;
  assign n31392 = ~n12861 & n31391;
  assign n31393 = ~n12240 & n31392;
  assign n31394 = ~n12973 & n31393;
  assign n31395 = n13109 & n31394;
  assign n31396 = n13095 & n31395;
  assign n31397 = n13134 & n31396;
  assign n31398 = ~n9717 & n26636;
  assign n31399 = ~n9913 & n31398;
  assign n31400 = n26634 & n31399;
  assign n31401 = ~n9929 & n31400;
  assign n31402 = ~n13824 & n31401;
  assign n31403 = ~n13823 & n31402;
  assign n31404 = ~n11266 & n31403;
  assign n31405 = ~n12861 & n31404;
  assign n31406 = ~n11588 & n31405;
  assign n31407 = ~n12973 & n31406;
  assign n31408 = n13054 & n31407;
  assign n31409 = n13095 & n31408;
  assign n31410 = n13858 & n31409;
  assign n31411 = ~n31397 & ~n31410;
  assign n31412 = pi071 & ~n2779;
  assign n31413 = ~n2780 & n31412;
  assign n31414 = ~n2778 & n31413;
  assign n31415 = ~n2543 & n31414;
  assign n31416 = n5772 & n31415;
  assign n31417 = ~n3066 & n31416;
  assign n31418 = ~n3983 & n31417;
  assign n31419 = ~n4003 & n31418;
  assign n31420 = ~n4024 & n31419;
  assign n31421 = ~n4999 & n31420;
  assign n31422 = ~n5827 & n31421;
  assign n31423 = ~n6893 & n31422;
  assign n31424 = ~n7890 & n31423;
  assign n31425 = ~n9131 & n31424;
  assign n31426 = ~n13144 & n31425;
  assign n31427 = ~n13143 & n31426;
  assign n31428 = ~n10278 & n31427;
  assign n31429 = ~n13142 & n31428;
  assign n31430 = ~n11662 & n31429;
  assign n31431 = ~n13141 & n31430;
  assign n31432 = n13165 & n31431;
  assign n31433 = n13140 & n31432;
  assign n31434 = n13190 & n31433;
  assign n31435 = pi119 & ~n5627;
  assign n31436 = n5687 & n31435;
  assign n31437 = n13580 & n31436;
  assign n31438 = ~n5808 & n31437;
  assign n31439 = ~n6056 & n31438;
  assign n31440 = ~n7073 & n31439;
  assign n31441 = ~n8179 & n31440;
  assign n31442 = ~n9344 & n31441;
  assign n31443 = ~n13517 & n31442;
  assign n31444 = ~n13516 & n31443;
  assign n31445 = ~n10594 & n31444;
  assign n31446 = ~n12861 & n31445;
  assign n31447 = ~n12005 & n31446;
  assign n31448 = ~n13515 & n31447;
  assign n31449 = n13532 & n31448;
  assign n31450 = n13514 & n31449;
  assign n31451 = n13557 & n31450;
  assign n31452 = ~n31434 & ~n31451;
  assign n31453 = n31411 & n31452;
  assign n31454 = n31381 & n31453;
  assign n31455 = n31308 & n31454;
  assign po120 = ~n31275 | ~n31455;
  assign n31457 = ~n11343 & n29206;
  assign n31458 = ~n12861 & n31457;
  assign n31459 = ~n11551 & n31458;
  assign n31460 = ~n12973 & n31459;
  assign n31461 = n13095 & n31460;
  assign n31462 = n13885 & n31461;
  assign n31463 = n13905 & n31462;
  assign n31464 = ~n10705 & n29215;
  assign n31465 = ~n12861 & n31464;
  assign n31466 = ~n12121 & n31465;
  assign n31467 = ~n13717 & n31466;
  assign n31468 = n13723 & n31467;
  assign n31469 = n13095 & n31468;
  assign n31470 = n13716 & n31469;
  assign n31471 = ~n31463 & ~n31470;
  assign n31472 = ~n11318 & n29129;
  assign n31473 = ~n12861 & n31472;
  assign n31474 = ~n12181 & n31473;
  assign n31475 = ~n13052 & n31474;
  assign n31476 = n13095 & n31475;
  assign n31477 = n13758 & n31476;
  assign n31478 = n13751 & n31477;
  assign n31479 = ~n10787 & n29107;
  assign n31480 = ~n12861 & n31479;
  assign n31481 = ~n11611 & n31480;
  assign n31482 = ~n12973 & n31481;
  assign n31483 = n13802 & n31482;
  assign n31484 = n13095 & n31483;
  assign n31485 = n13819 & n31484;
  assign n31486 = ~n31478 & ~n31485;
  assign n31487 = n31471 & n31486;
  assign n31488 = n13731 & n24849;
  assign n31489 = ~n7869 & n31488;
  assign n31490 = ~n8346 & n31489;
  assign n31491 = ~n9485 & n31490;
  assign n31492 = ~n13653 & n31491;
  assign n31493 = ~n13652 & n31492;
  assign n31494 = ~n10741 & n31493;
  assign n31495 = ~n12861 & n31494;
  assign n31496 = ~n12158 & n31495;
  assign n31497 = ~n13052 & n31496;
  assign n31498 = n13667 & n31497;
  assign n31499 = n13095 & n31498;
  assign n31500 = n13692 & n31499;
  assign n31501 = ~n12041 & n29047;
  assign n31502 = ~n12861 & n31501;
  assign n31503 = n13094 & n31502;
  assign n31504 = n13577 & n31503;
  assign n31505 = n13572 & n31504;
  assign n31506 = ~n13312 & n28978;
  assign n31507 = ~n13310 & n31506;
  assign n31508 = n13317 & n31507;
  assign n31509 = pi232 & ~n501;
  assign n31510 = n14255 & n31509;
  assign n31511 = n14253 & n31510;
  assign n31512 = n31154 & n31511;
  assign n31513 = n31162 & n31512;
  assign n31514 = ~n1172 & n31513;
  assign n31515 = ~n996 & n31514;
  assign n31516 = ~n2306 & n31515;
  assign n31517 = n3819 & n31516;
  assign n31518 = n14139 & n31517;
  assign n31519 = n12583 & n31518;
  assign n31520 = n14252 & n31519;
  assign n31521 = n14242 & n31520;
  assign n31522 = n14431 & n31521;
  assign n31523 = ~n7236 & n31522;
  assign n31524 = ~n6137 & n31523;
  assign n31525 = n6193 & n31524;
  assign n31526 = n6134 & n31525;
  assign n31527 = ~n8867 & n31526;
  assign n31528 = ~n7235 & n31527;
  assign n31529 = n7296 & n31528;
  assign n31530 = n7231 & n31529;
  assign n31531 = ~n10027 & n31530;
  assign n31532 = ~n8866 & n31531;
  assign n31533 = n8898 & n31532;
  assign n31534 = n8863 & n31533;
  assign n31535 = pi240 & ~n501;
  assign n31536 = n14188 & n31535;
  assign n31537 = n31189 & n31536;
  assign n31538 = n31196 & n31537;
  assign n31539 = ~n1172 & n31538;
  assign n31540 = ~n996 & n31539;
  assign n31541 = ~n2306 & n31540;
  assign n31542 = n3819 & n31541;
  assign n31543 = n3821 & n31542;
  assign n31544 = n14186 & n31543;
  assign n31545 = n14229 & n31544;
  assign n31546 = n14184 & n31545;
  assign n31547 = n14180 & n31546;
  assign n31548 = ~n7236 & n31547;
  assign n31549 = ~n6137 & n31548;
  assign n31550 = n6193 & n31549;
  assign n31551 = n6134 & n31550;
  assign n31552 = ~n8867 & n31551;
  assign n31553 = ~n7235 & n31552;
  assign n31554 = n7296 & n31553;
  assign n31555 = n7231 & n31554;
  assign n31556 = ~n10027 & n31555;
  assign n31557 = ~n8866 & n31556;
  assign n31558 = n8898 & n31557;
  assign n31559 = n8863 & n31558;
  assign n31560 = ~n31534 & ~n31559;
  assign n31561 = ~n10788 & ~n31560;
  assign n31562 = ~n10026 & n31561;
  assign n31563 = n10072 & n31562;
  assign n31564 = n10021 & n31563;
  assign n31565 = ~n31508 & ~n31564;
  assign n31566 = ~n31505 & n31565;
  assign n31567 = ~n11860 & n28974;
  assign n31568 = ~n12861 & n31567;
  assign n31569 = ~n13399 & n31568;
  assign n31570 = n13406 & n31569;
  assign n31571 = ~n11959 & n29042;
  assign n31572 = ~n12861 & n31571;
  assign n31573 = ~n12950 & n31572;
  assign n31574 = n13491 & n31573;
  assign n31575 = n13486 & n31574;
  assign n31576 = ~n31570 & ~n31575;
  assign n31577 = n31566 & n31576;
  assign n31578 = ~n31500 & n31577;
  assign n31579 = pi184 & ~n9717;
  assign n31580 = ~n9913 & n31579;
  assign n31581 = n9856 & n31580;
  assign n31582 = ~n9929 & n31581;
  assign n31583 = ~n13824 & n31582;
  assign n31584 = ~n13823 & n31583;
  assign n31585 = ~n11266 & n31584;
  assign n31586 = ~n12861 & n31585;
  assign n31587 = ~n11588 & n31586;
  assign n31588 = ~n12973 & n31587;
  assign n31589 = n13054 & n31588;
  assign n31590 = n13095 & n31589;
  assign n31591 = n13858 & n31590;
  assign n31592 = pi168 & ~n8574;
  assign n31593 = n11377 & n31592;
  assign n31594 = n9942 & n31593;
  assign n31595 = ~n8834 & n31594;
  assign n31596 = ~n10002 & n31595;
  assign n31597 = ~n13097 & n31596;
  assign n31598 = ~n13096 & n31597;
  assign n31599 = ~n11297 & n31598;
  assign n31600 = ~n12861 & n31599;
  assign n31601 = ~n12240 & n31600;
  assign n31602 = ~n12973 & n31601;
  assign n31603 = n13109 & n31602;
  assign n31604 = n13095 & n31603;
  assign n31605 = n13134 & n31604;
  assign n31606 = ~n31591 & ~n31605;
  assign n31607 = n31578 & n31606;
  assign n31608 = n31487 & n31607;
  assign n31609 = pi216 & ~n12671;
  assign n31610 = ~n12811 & n31609;
  assign n31611 = n13912 & n31610;
  assign n31612 = ~n12902 & n31611;
  assign n31613 = ~n13908 & n31612;
  assign n31614 = ~n12861 & n31613;
  assign n31615 = ~n12860 & n31614;
  assign n31616 = n12952 & n31615;
  assign n31617 = n13919 & n31616;
  assign n31618 = n14008 & n31617;
  assign n31619 = n7175 & n27007;
  assign n31620 = n13694 & n31619;
  assign n31621 = ~n6784 & n31620;
  assign n31622 = ~n7158 & n31621;
  assign n31623 = ~n8250 & n31622;
  assign n31624 = ~n9414 & n31623;
  assign n31625 = ~n13602 & n31624;
  assign n31626 = ~n13601 & n31625;
  assign n31627 = ~n10667 & n31626;
  assign n31628 = ~n12861 & n31627;
  assign n31629 = ~n12083 & n31628;
  assign n31630 = ~n13600 & n31629;
  assign n31631 = n13618 & n31630;
  assign n31632 = n13095 & n31631;
  assign n31633 = n13643 & n31632;
  assign n31634 = n13408 & n26788;
  assign n31635 = ~n3940 & n31634;
  assign n31636 = ~n4001 & n31635;
  assign n31637 = ~n5043 & n31636;
  assign n31638 = ~n5943 & n31637;
  assign n31639 = ~n6951 & n31638;
  assign n31640 = ~n8037 & n31639;
  assign n31641 = ~n9200 & n31640;
  assign n31642 = ~n13348 & n31641;
  assign n31643 = ~n13347 & n31642;
  assign n31644 = ~n10445 & n31643;
  assign n31645 = ~n12861 & n31644;
  assign n31646 = ~n11846 & n31645;
  assign n31647 = ~n13346 & n31646;
  assign n31648 = n13367 & n31647;
  assign n31649 = n13345 & n31648;
  assign n31650 = n13392 & n31649;
  assign n31651 = ~n31633 & ~n31650;
  assign n31652 = ~n31618 & n31651;
  assign n31653 = pi056 & ~n1679;
  assign n31654 = n1741 & n31653;
  assign n31655 = n13259 & n31654;
  assign n31656 = ~n2242 & n31655;
  assign n31657 = ~n3095 & n31656;
  assign n31658 = ~n3997 & n31657;
  assign n31659 = ~n4003 & n31658;
  assign n31660 = ~n4837 & n31659;
  assign n31661 = ~n5822 & n31660;
  assign n31662 = ~n6820 & n31661;
  assign n31663 = ~n7785 & n31662;
  assign n31664 = ~n9027 & n31663;
  assign n31665 = ~n10245 & n31664;
  assign n31666 = ~n13258 & n31665;
  assign n31667 = ~n13257 & n31666;
  assign n31668 = ~n11536 & n31667;
  assign n31669 = ~n13256 & n31668;
  assign n31670 = ~n13036 & n31669;
  assign n31671 = ~n13255 & n31670;
  assign n31672 = n13281 & n31671;
  assign n31673 = n13254 & n31672;
  assign n31674 = n13306 & n31673;
  assign n31675 = pi224 & ~n12946;
  assign n31676 = ~n12903 & n31675;
  assign n31677 = ~n12861 & n31676;
  assign n31678 = ~n12860 & n31677;
  assign n31679 = n12952 & n31678;
  assign n31680 = n12975 & n31679;
  assign n31681 = n13092 & n31680;
  assign n31682 = ~n31674 & ~n31681;
  assign n31683 = n13319 & n24860;
  assign n31684 = ~n3066 & n31683;
  assign n31685 = ~n3983 & n31684;
  assign n31686 = ~n4003 & n31685;
  assign n31687 = ~n4024 & n31686;
  assign n31688 = ~n4999 & n31687;
  assign n31689 = ~n5827 & n31688;
  assign n31690 = ~n6893 & n31689;
  assign n31691 = ~n7890 & n31690;
  assign n31692 = ~n9131 & n31691;
  assign n31693 = ~n13144 & n31692;
  assign n31694 = ~n13143 & n31693;
  assign n31695 = ~n10278 & n31694;
  assign n31696 = ~n13142 & n31695;
  assign n31697 = ~n11662 & n31696;
  assign n31698 = ~n13141 & n31697;
  assign n31699 = n13165 & n31698;
  assign n31700 = n13140 & n31699;
  assign n31701 = n13190 & n31700;
  assign n31702 = n13494 & n26816;
  assign n31703 = ~n4817 & n31702;
  assign n31704 = ~n4902 & n31703;
  assign n31705 = ~n6001 & n31704;
  assign n31706 = ~n7014 & n31705;
  assign n31707 = ~n8114 & n31706;
  assign n31708 = ~n9276 & n31707;
  assign n31709 = ~n13438 & n31708;
  assign n31710 = ~n13437 & n31709;
  assign n31711 = ~n10523 & n31710;
  assign n31712 = ~n12861 & n31711;
  assign n31713 = ~n11928 & n31712;
  assign n31714 = ~n13436 & n31713;
  assign n31715 = n13453 & n31714;
  assign n31716 = n13435 & n31715;
  assign n31717 = n13478 & n31716;
  assign n31718 = ~n31701 & ~n31717;
  assign n31719 = n31682 & n31718;
  assign n31720 = pi200 & ~n10909;
  assign n31721 = ~n11168 & n31720;
  assign n31722 = n11135 & n31721;
  assign n31723 = ~n11188 & n31722;
  assign n31724 = ~n14011 & n31723;
  assign n31725 = ~n14010 & n31724;
  assign n31726 = ~n12861 & n31725;
  assign n31727 = ~n12380 & n31726;
  assign n31728 = ~n12972 & n31727;
  assign n31729 = n14020 & n31728;
  assign n31730 = n13095 & n31729;
  assign n31731 = n14044 & n31730;
  assign n31732 = n13202 & n26953;
  assign n31733 = ~n1372 & n31732;
  assign n31734 = ~n2243 & n31733;
  assign n31735 = ~n3104 & n31734;
  assign n31736 = ~n3971 & n31735;
  assign n31737 = ~n4003 & n31736;
  assign n31738 = ~n4872 & n31737;
  assign n31739 = ~n5801 & n31738;
  assign n31740 = ~n6739 & n31739;
  assign n31741 = ~n7807 & n31740;
  assign n31742 = ~n8989 & n31741;
  assign n31743 = ~n10273 & n31742;
  assign n31744 = ~n13200 & n31743;
  assign n31745 = ~n13199 & n31744;
  assign n31746 = ~n11499 & n31745;
  assign n31747 = ~n13198 & n31746;
  assign n31748 = ~n13076 & n31747;
  assign n31749 = ~n13197 & n31748;
  assign n31750 = n13223 & n31749;
  assign n31751 = n13196 & n31750;
  assign n31752 = n13248 & n31751;
  assign n31753 = ~n31731 & ~n31752;
  assign n31754 = ~n12861 & n29169;
  assign n31755 = ~n12471 & n31754;
  assign n31756 = ~n12972 & n31755;
  assign n31757 = n14020 & n31756;
  assign n31758 = n13095 & n31757;
  assign n31759 = n14072 & n31758;
  assign n31760 = pi120 & ~n5627;
  assign n31761 = n5687 & n31760;
  assign n31762 = n13580 & n31761;
  assign n31763 = ~n5808 & n31762;
  assign n31764 = ~n6056 & n31763;
  assign n31765 = ~n7073 & n31764;
  assign n31766 = ~n8179 & n31765;
  assign n31767 = ~n9344 & n31766;
  assign n31768 = ~n13517 & n31767;
  assign n31769 = ~n13516 & n31768;
  assign n31770 = ~n10594 & n31769;
  assign n31771 = ~n12861 & n31770;
  assign n31772 = ~n12005 & n31771;
  assign n31773 = ~n13515 & n31772;
  assign n31774 = n13532 & n31773;
  assign n31775 = n13514 & n31774;
  assign n31776 = n13557 & n31775;
  assign n31777 = ~n31759 & ~n31776;
  assign n31778 = n31753 & n31777;
  assign n31779 = n31719 & n31778;
  assign n31780 = n31652 & n31779;
  assign po121 = ~n31608 | ~n31780;
  assign n31782 = ~n10787 & n29481;
  assign n31783 = ~n12861 & n31782;
  assign n31784 = ~n11611 & n31783;
  assign n31785 = ~n12973 & n31784;
  assign n31786 = n13802 & n31785;
  assign n31787 = n13095 & n31786;
  assign n31788 = n13819 & n31787;
  assign n31789 = ~n10705 & n29550;
  assign n31790 = ~n12861 & n31789;
  assign n31791 = ~n12121 & n31790;
  assign n31792 = ~n13717 & n31791;
  assign n31793 = n13723 & n31792;
  assign n31794 = n13095 & n31793;
  assign n31795 = n13716 & n31794;
  assign n31796 = ~n31788 & ~n31795;
  assign n31797 = ~n11318 & n29355;
  assign n31798 = ~n12861 & n31797;
  assign n31799 = ~n12181 & n31798;
  assign n31800 = ~n13052 & n31799;
  assign n31801 = n13095 & n31800;
  assign n31802 = n13758 & n31801;
  assign n31803 = n13751 & n31802;
  assign n31804 = ~n11343 & n29518;
  assign n31805 = ~n12861 & n31804;
  assign n31806 = ~n11551 & n31805;
  assign n31807 = ~n12973 & n31806;
  assign n31808 = n13095 & n31807;
  assign n31809 = n13885 & n31808;
  assign n31810 = n13905 & n31809;
  assign n31811 = ~n31803 & ~n31810;
  assign n31812 = n31796 & n31811;
  assign n31813 = pi057 & ~n1679;
  assign n31814 = n1741 & n31813;
  assign n31815 = n13259 & n31814;
  assign n31816 = ~n2242 & n31815;
  assign n31817 = ~n3095 & n31816;
  assign n31818 = ~n3997 & n31817;
  assign n31819 = ~n4003 & n31818;
  assign n31820 = ~n4837 & n31819;
  assign n31821 = ~n5822 & n31820;
  assign n31822 = ~n6820 & n31821;
  assign n31823 = ~n7785 & n31822;
  assign n31824 = ~n9027 & n31823;
  assign n31825 = ~n10245 & n31824;
  assign n31826 = ~n13258 & n31825;
  assign n31827 = ~n13257 & n31826;
  assign n31828 = ~n11536 & n31827;
  assign n31829 = ~n13256 & n31828;
  assign n31830 = ~n13036 & n31829;
  assign n31831 = ~n13255 & n31830;
  assign n31832 = n13281 & n31831;
  assign n31833 = n13254 & n31832;
  assign n31834 = n13306 & n31833;
  assign n31835 = ~n11860 & n29275;
  assign n31836 = ~n12861 & n31835;
  assign n31837 = ~n13399 & n31836;
  assign n31838 = n13406 & n31837;
  assign n31839 = ~n13312 & n29279;
  assign n31840 = ~n13310 & n31839;
  assign n31841 = n13317 & n31840;
  assign n31842 = pi241 & ~n501;
  assign n31843 = n14188 & n31842;
  assign n31844 = n31189 & n31843;
  assign n31845 = n31196 & n31844;
  assign n31846 = ~n1172 & n31845;
  assign n31847 = ~n996 & n31846;
  assign n31848 = ~n2306 & n31847;
  assign n31849 = n3819 & n31848;
  assign n31850 = n3821 & n31849;
  assign n31851 = n14186 & n31850;
  assign n31852 = n14229 & n31851;
  assign n31853 = n14184 & n31852;
  assign n31854 = n14180 & n31853;
  assign n31855 = ~n7236 & n31854;
  assign n31856 = ~n6137 & n31855;
  assign n31857 = n6193 & n31856;
  assign n31858 = n6134 & n31857;
  assign n31859 = ~n8867 & n31858;
  assign n31860 = ~n7235 & n31859;
  assign n31861 = n7296 & n31860;
  assign n31862 = n7231 & n31861;
  assign n31863 = ~n10027 & n31862;
  assign n31864 = ~n8866 & n31863;
  assign n31865 = n8898 & n31864;
  assign n31866 = n8863 & n31865;
  assign n31867 = pi233 & ~n501;
  assign n31868 = n14255 & n31867;
  assign n31869 = n14253 & n31868;
  assign n31870 = n31154 & n31869;
  assign n31871 = n31162 & n31870;
  assign n31872 = ~n1172 & n31871;
  assign n31873 = ~n996 & n31872;
  assign n31874 = ~n2306 & n31873;
  assign n31875 = n3819 & n31874;
  assign n31876 = n14139 & n31875;
  assign n31877 = n12583 & n31876;
  assign n31878 = n14252 & n31877;
  assign n31879 = n14242 & n31878;
  assign n31880 = n14431 & n31879;
  assign n31881 = ~n7236 & n31880;
  assign n31882 = ~n6137 & n31881;
  assign n31883 = n6193 & n31882;
  assign n31884 = n6134 & n31883;
  assign n31885 = ~n8867 & n31884;
  assign n31886 = ~n7235 & n31885;
  assign n31887 = n7296 & n31886;
  assign n31888 = n7231 & n31887;
  assign n31889 = ~n10027 & n31888;
  assign n31890 = ~n8866 & n31889;
  assign n31891 = n8898 & n31890;
  assign n31892 = n8863 & n31891;
  assign n31893 = ~n31866 & ~n31892;
  assign n31894 = ~n10788 & ~n31893;
  assign n31895 = ~n10026 & n31894;
  assign n31896 = n10072 & n31895;
  assign n31897 = n10021 & n31896;
  assign n31898 = ~n31841 & ~n31897;
  assign n31899 = ~n31838 & n31898;
  assign n31900 = ~n11959 & n29343;
  assign n31901 = ~n12861 & n31900;
  assign n31902 = ~n12950 & n31901;
  assign n31903 = n13491 & n31902;
  assign n31904 = n13486 & n31903;
  assign n31905 = ~n12041 & n29348;
  assign n31906 = ~n12861 & n31905;
  assign n31907 = n13094 & n31906;
  assign n31908 = n13577 & n31907;
  assign n31909 = n13572 & n31908;
  assign n31910 = ~n31904 & ~n31909;
  assign n31911 = n31899 & n31910;
  assign n31912 = ~n31834 & n31911;
  assign n31913 = n13731 & n25226;
  assign n31914 = ~n7869 & n31913;
  assign n31915 = ~n8346 & n31914;
  assign n31916 = ~n9485 & n31915;
  assign n31917 = ~n13653 & n31916;
  assign n31918 = ~n13652 & n31917;
  assign n31919 = ~n10741 & n31918;
  assign n31920 = ~n12861 & n31919;
  assign n31921 = ~n12158 & n31920;
  assign n31922 = ~n13052 & n31921;
  assign n31923 = n13667 & n31922;
  assign n31924 = n13095 & n31923;
  assign n31925 = n13692 & n31924;
  assign n31926 = n13202 & n27216;
  assign n31927 = ~n1372 & n31926;
  assign n31928 = ~n2243 & n31927;
  assign n31929 = ~n3104 & n31928;
  assign n31930 = ~n3971 & n31929;
  assign n31931 = ~n4003 & n31930;
  assign n31932 = ~n4872 & n31931;
  assign n31933 = ~n5801 & n31932;
  assign n31934 = ~n6739 & n31933;
  assign n31935 = ~n7807 & n31934;
  assign n31936 = ~n8989 & n31935;
  assign n31937 = ~n10273 & n31936;
  assign n31938 = ~n13200 & n31937;
  assign n31939 = ~n13199 & n31938;
  assign n31940 = ~n11499 & n31939;
  assign n31941 = ~n13198 & n31940;
  assign n31942 = ~n13076 & n31941;
  assign n31943 = ~n13197 & n31942;
  assign n31944 = n13223 & n31943;
  assign n31945 = n13196 & n31944;
  assign n31946 = n13248 & n31945;
  assign n31947 = ~n31925 & ~n31946;
  assign n31948 = n31912 & n31947;
  assign n31949 = n31812 & n31948;
  assign n31950 = n7175 & n27238;
  assign n31951 = n13694 & n31950;
  assign n31952 = ~n6784 & n31951;
  assign n31953 = ~n7158 & n31952;
  assign n31954 = ~n8250 & n31953;
  assign n31955 = ~n9414 & n31954;
  assign n31956 = ~n13602 & n31955;
  assign n31957 = ~n13601 & n31956;
  assign n31958 = ~n10667 & n31957;
  assign n31959 = ~n12861 & n31958;
  assign n31960 = ~n12083 & n31959;
  assign n31961 = ~n13600 & n31960;
  assign n31962 = n13618 & n31961;
  assign n31963 = n13095 & n31962;
  assign n31964 = n13643 & n31963;
  assign n31965 = n13319 & n25206;
  assign n31966 = ~n3066 & n31965;
  assign n31967 = ~n3983 & n31966;
  assign n31968 = ~n4003 & n31967;
  assign n31969 = ~n4024 & n31968;
  assign n31970 = ~n4999 & n31969;
  assign n31971 = ~n5827 & n31970;
  assign n31972 = ~n6893 & n31971;
  assign n31973 = ~n7890 & n31972;
  assign n31974 = ~n9131 & n31973;
  assign n31975 = ~n13144 & n31974;
  assign n31976 = ~n13143 & n31975;
  assign n31977 = ~n10278 & n31976;
  assign n31978 = ~n13142 & n31977;
  assign n31979 = ~n11662 & n31978;
  assign n31980 = ~n13141 & n31979;
  assign n31981 = n13165 & n31980;
  assign n31982 = n13140 & n31981;
  assign n31983 = n13190 & n31982;
  assign n31984 = pi121 & ~n5627;
  assign n31985 = n5687 & n31984;
  assign n31986 = n13580 & n31985;
  assign n31987 = ~n5808 & n31986;
  assign n31988 = ~n6056 & n31987;
  assign n31989 = ~n7073 & n31988;
  assign n31990 = ~n8179 & n31989;
  assign n31991 = ~n9344 & n31990;
  assign n31992 = ~n13517 & n31991;
  assign n31993 = ~n13516 & n31992;
  assign n31994 = ~n10594 & n31993;
  assign n31995 = ~n12861 & n31994;
  assign n31996 = ~n12005 & n31995;
  assign n31997 = ~n13515 & n31996;
  assign n31998 = n13532 & n31997;
  assign n31999 = n13514 & n31998;
  assign n32000 = n13557 & n31999;
  assign n32001 = ~n31983 & ~n32000;
  assign n32002 = ~n31964 & n32001;
  assign n32003 = pi169 & ~n8574;
  assign n32004 = n11377 & n32003;
  assign n32005 = n9942 & n32004;
  assign n32006 = ~n8834 & n32005;
  assign n32007 = ~n10002 & n32006;
  assign n32008 = ~n13097 & n32007;
  assign n32009 = ~n13096 & n32008;
  assign n32010 = ~n11297 & n32009;
  assign n32011 = ~n12861 & n32010;
  assign n32012 = ~n12240 & n32011;
  assign n32013 = ~n12973 & n32012;
  assign n32014 = n13109 & n32013;
  assign n32015 = n13095 & n32014;
  assign n32016 = n13134 & n32015;
  assign n32017 = pi225 & ~n12946;
  assign n32018 = ~n12903 & n32017;
  assign n32019 = ~n12861 & n32018;
  assign n32020 = ~n12860 & n32019;
  assign n32021 = n12952 & n32020;
  assign n32022 = n12975 & n32021;
  assign n32023 = n13092 & n32022;
  assign n32024 = ~n32016 & ~n32023;
  assign n32025 = pi217 & ~n12671;
  assign n32026 = ~n12811 & n32025;
  assign n32027 = n13912 & n32026;
  assign n32028 = ~n12902 & n32027;
  assign n32029 = ~n13908 & n32028;
  assign n32030 = ~n12861 & n32029;
  assign n32031 = ~n12860 & n32030;
  assign n32032 = n12952 & n32031;
  assign n32033 = n13919 & n32032;
  assign n32034 = n14008 & n32033;
  assign n32035 = ~n12861 & n29527;
  assign n32036 = ~n12471 & n32035;
  assign n32037 = ~n12972 & n32036;
  assign n32038 = n14020 & n32037;
  assign n32039 = n13095 & n32038;
  assign n32040 = n14072 & n32039;
  assign n32041 = ~n32034 & ~n32040;
  assign n32042 = n32024 & n32041;
  assign n32043 = pi201 & ~n10909;
  assign n32044 = ~n11168 & n32043;
  assign n32045 = n11135 & n32044;
  assign n32046 = ~n11188 & n32045;
  assign n32047 = ~n14011 & n32046;
  assign n32048 = ~n14010 & n32047;
  assign n32049 = ~n12861 & n32048;
  assign n32050 = ~n12380 & n32049;
  assign n32051 = ~n12972 & n32050;
  assign n32052 = n14020 & n32051;
  assign n32053 = n13095 & n32052;
  assign n32054 = n14044 & n32053;
  assign n32055 = n13408 & n27271;
  assign n32056 = ~n3940 & n32055;
  assign n32057 = ~n4001 & n32056;
  assign n32058 = ~n5043 & n32057;
  assign n32059 = ~n5943 & n32058;
  assign n32060 = ~n6951 & n32059;
  assign n32061 = ~n8037 & n32060;
  assign n32062 = ~n9200 & n32061;
  assign n32063 = ~n13348 & n32062;
  assign n32064 = ~n13347 & n32063;
  assign n32065 = ~n10445 & n32064;
  assign n32066 = ~n12861 & n32065;
  assign n32067 = ~n11846 & n32066;
  assign n32068 = ~n13346 & n32067;
  assign n32069 = n13367 & n32068;
  assign n32070 = n13345 & n32069;
  assign n32071 = n13392 & n32070;
  assign n32072 = ~n32054 & ~n32071;
  assign n32073 = pi185 & ~n9717;
  assign n32074 = ~n9913 & n32073;
  assign n32075 = n9856 & n32074;
  assign n32076 = ~n9929 & n32075;
  assign n32077 = ~n13824 & n32076;
  assign n32078 = ~n13823 & n32077;
  assign n32079 = ~n11266 & n32078;
  assign n32080 = ~n12861 & n32079;
  assign n32081 = ~n11588 & n32080;
  assign n32082 = ~n12973 & n32081;
  assign n32083 = n13054 & n32082;
  assign n32084 = n13095 & n32083;
  assign n32085 = n13858 & n32084;
  assign n32086 = n13494 & n27054;
  assign n32087 = ~n4817 & n32086;
  assign n32088 = ~n4902 & n32087;
  assign n32089 = ~n6001 & n32088;
  assign n32090 = ~n7014 & n32089;
  assign n32091 = ~n8114 & n32090;
  assign n32092 = ~n9276 & n32091;
  assign n32093 = ~n13438 & n32092;
  assign n32094 = ~n13437 & n32093;
  assign n32095 = ~n10523 & n32094;
  assign n32096 = ~n12861 & n32095;
  assign n32097 = ~n11928 & n32096;
  assign n32098 = ~n13436 & n32097;
  assign n32099 = n13453 & n32098;
  assign n32100 = n13435 & n32099;
  assign n32101 = n13478 & n32100;
  assign n32102 = ~n32085 & ~n32101;
  assign n32103 = n32072 & n32102;
  assign n32104 = n32042 & n32103;
  assign n32105 = n32002 & n32104;
  assign po122 = ~n31949 | ~n32105;
  assign n32107 = ~n10787 & n29828;
  assign n32108 = ~n12861 & n32107;
  assign n32109 = ~n11611 & n32108;
  assign n32110 = ~n12973 & n32109;
  assign n32111 = n13802 & n32110;
  assign n32112 = n13095 & n32111;
  assign n32113 = n13819 & n32112;
  assign n32114 = ~n10705 & n29711;
  assign n32115 = ~n12861 & n32114;
  assign n32116 = ~n12121 & n32115;
  assign n32117 = ~n13717 & n32116;
  assign n32118 = n13723 & n32117;
  assign n32119 = n13095 & n32118;
  assign n32120 = n13716 & n32119;
  assign n32121 = ~n32113 & ~n32120;
  assign n32122 = ~n11318 & n29782;
  assign n32123 = ~n12861 & n32122;
  assign n32124 = ~n12181 & n32123;
  assign n32125 = ~n13052 & n32124;
  assign n32126 = n13095 & n32125;
  assign n32127 = n13758 & n32126;
  assign n32128 = n13751 & n32127;
  assign n32129 = ~n11343 & n29802;
  assign n32130 = ~n12861 & n32129;
  assign n32131 = ~n11551 & n32130;
  assign n32132 = ~n12973 & n32131;
  assign n32133 = n13095 & n32132;
  assign n32134 = n13885 & n32133;
  assign n32135 = n13905 & n32134;
  assign n32136 = ~n32128 & ~n32135;
  assign n32137 = n32121 & n32136;
  assign n32138 = n13731 & n25457;
  assign n32139 = ~n7869 & n32138;
  assign n32140 = ~n8346 & n32139;
  assign n32141 = ~n9485 & n32140;
  assign n32142 = ~n13653 & n32141;
  assign n32143 = ~n13652 & n32142;
  assign n32144 = ~n10741 & n32143;
  assign n32145 = ~n12861 & n32144;
  assign n32146 = ~n12158 & n32145;
  assign n32147 = ~n13052 & n32146;
  assign n32148 = n13667 & n32147;
  assign n32149 = n13095 & n32148;
  assign n32150 = n13692 & n32149;
  assign n32151 = ~n11860 & n29576;
  assign n32152 = ~n12861 & n32151;
  assign n32153 = ~n13399 & n32152;
  assign n32154 = n13406 & n32153;
  assign n32155 = ~n13312 & n29580;
  assign n32156 = ~n13310 & n32155;
  assign n32157 = n13317 & n32156;
  assign n32158 = pi234 & ~n501;
  assign n32159 = n14255 & n32158;
  assign n32160 = n14253 & n32159;
  assign n32161 = n31154 & n32160;
  assign n32162 = n31162 & n32161;
  assign n32163 = ~n1172 & n32162;
  assign n32164 = ~n996 & n32163;
  assign n32165 = ~n2306 & n32164;
  assign n32166 = n3819 & n32165;
  assign n32167 = n14139 & n32166;
  assign n32168 = n12583 & n32167;
  assign n32169 = n14252 & n32168;
  assign n32170 = n14242 & n32169;
  assign n32171 = n14431 & n32170;
  assign n32172 = ~n7236 & n32171;
  assign n32173 = ~n6137 & n32172;
  assign n32174 = n6193 & n32173;
  assign n32175 = n6134 & n32174;
  assign n32176 = ~n8867 & n32175;
  assign n32177 = ~n7235 & n32176;
  assign n32178 = n7296 & n32177;
  assign n32179 = n7231 & n32178;
  assign n32180 = ~n10027 & n32179;
  assign n32181 = ~n8866 & n32180;
  assign n32182 = n8898 & n32181;
  assign n32183 = n8863 & n32182;
  assign n32184 = pi242 & ~n501;
  assign n32185 = n14188 & n32184;
  assign n32186 = n31189 & n32185;
  assign n32187 = n31196 & n32186;
  assign n32188 = ~n1172 & n32187;
  assign n32189 = ~n996 & n32188;
  assign n32190 = ~n2306 & n32189;
  assign n32191 = n3819 & n32190;
  assign n32192 = n3821 & n32191;
  assign n32193 = n14186 & n32192;
  assign n32194 = n14229 & n32193;
  assign n32195 = n14184 & n32194;
  assign n32196 = n14180 & n32195;
  assign n32197 = ~n7236 & n32196;
  assign n32198 = ~n6137 & n32197;
  assign n32199 = n6193 & n32198;
  assign n32200 = n6134 & n32199;
  assign n32201 = ~n8867 & n32200;
  assign n32202 = ~n7235 & n32201;
  assign n32203 = n7296 & n32202;
  assign n32204 = n7231 & n32203;
  assign n32205 = ~n10027 & n32204;
  assign n32206 = ~n8866 & n32205;
  assign n32207 = n8898 & n32206;
  assign n32208 = n8863 & n32207;
  assign n32209 = ~n32183 & ~n32208;
  assign n32210 = ~n10788 & ~n32209;
  assign n32211 = ~n10026 & n32210;
  assign n32212 = n10072 & n32211;
  assign n32213 = n10021 & n32212;
  assign n32214 = ~n32157 & ~n32213;
  assign n32215 = ~n32154 & n32214;
  assign n32216 = ~n11959 & n29644;
  assign n32217 = ~n12861 & n32216;
  assign n32218 = ~n12950 & n32217;
  assign n32219 = n13491 & n32218;
  assign n32220 = n13486 & n32219;
  assign n32221 = ~n12041 & n29649;
  assign n32222 = ~n12861 & n32221;
  assign n32223 = n13094 & n32222;
  assign n32224 = n13577 & n32223;
  assign n32225 = n13572 & n32224;
  assign n32226 = ~n32220 & ~n32225;
  assign n32227 = n32215 & n32226;
  assign n32228 = ~n32150 & n32227;
  assign n32229 = pi058 & ~n1679;
  assign n32230 = n1741 & n32229;
  assign n32231 = n13259 & n32230;
  assign n32232 = ~n2242 & n32231;
  assign n32233 = ~n3095 & n32232;
  assign n32234 = ~n3997 & n32233;
  assign n32235 = ~n4003 & n32234;
  assign n32236 = ~n4837 & n32235;
  assign n32237 = ~n5822 & n32236;
  assign n32238 = ~n6820 & n32237;
  assign n32239 = ~n7785 & n32238;
  assign n32240 = ~n9027 & n32239;
  assign n32241 = ~n10245 & n32240;
  assign n32242 = ~n13258 & n32241;
  assign n32243 = ~n13257 & n32242;
  assign n32244 = ~n11536 & n32243;
  assign n32245 = ~n13256 & n32244;
  assign n32246 = ~n13036 & n32245;
  assign n32247 = ~n13255 & n32246;
  assign n32248 = n13281 & n32247;
  assign n32249 = n13254 & n32248;
  assign n32250 = n13306 & n32249;
  assign n32251 = n13202 & n27478;
  assign n32252 = ~n1372 & n32251;
  assign n32253 = ~n2243 & n32252;
  assign n32254 = ~n3104 & n32253;
  assign n32255 = ~n3971 & n32254;
  assign n32256 = ~n4003 & n32255;
  assign n32257 = ~n4872 & n32256;
  assign n32258 = ~n5801 & n32257;
  assign n32259 = ~n6739 & n32258;
  assign n32260 = ~n7807 & n32259;
  assign n32261 = ~n8989 & n32260;
  assign n32262 = ~n10273 & n32261;
  assign n32263 = ~n13200 & n32262;
  assign n32264 = ~n13199 & n32263;
  assign n32265 = ~n11499 & n32264;
  assign n32266 = ~n13198 & n32265;
  assign n32267 = ~n13076 & n32266;
  assign n32268 = ~n13197 & n32267;
  assign n32269 = n13223 & n32268;
  assign n32270 = n13196 & n32269;
  assign n32271 = n13248 & n32270;
  assign n32272 = ~n32250 & ~n32271;
  assign n32273 = n32228 & n32272;
  assign n32274 = n32137 & n32273;
  assign n32275 = n7175 & n27435;
  assign n32276 = n13694 & n32275;
  assign n32277 = ~n6784 & n32276;
  assign n32278 = ~n7158 & n32277;
  assign n32279 = ~n8250 & n32278;
  assign n32280 = ~n9414 & n32279;
  assign n32281 = ~n13602 & n32280;
  assign n32282 = ~n13601 & n32281;
  assign n32283 = ~n10667 & n32282;
  assign n32284 = ~n12861 & n32283;
  assign n32285 = ~n12083 & n32284;
  assign n32286 = ~n13600 & n32285;
  assign n32287 = n13618 & n32286;
  assign n32288 = n13095 & n32287;
  assign n32289 = n13643 & n32288;
  assign n32290 = n13494 & n27538;
  assign n32291 = ~n4817 & n32290;
  assign n32292 = ~n4902 & n32291;
  assign n32293 = ~n6001 & n32292;
  assign n32294 = ~n7014 & n32293;
  assign n32295 = ~n8114 & n32294;
  assign n32296 = ~n9276 & n32295;
  assign n32297 = ~n13438 & n32296;
  assign n32298 = ~n13437 & n32297;
  assign n32299 = ~n10523 & n32298;
  assign n32300 = ~n12861 & n32299;
  assign n32301 = ~n11928 & n32300;
  assign n32302 = ~n13436 & n32301;
  assign n32303 = n13453 & n32302;
  assign n32304 = n13435 & n32303;
  assign n32305 = n13478 & n32304;
  assign n32306 = pi122 & ~n5627;
  assign n32307 = n5687 & n32306;
  assign n32308 = n13580 & n32307;
  assign n32309 = ~n5808 & n32308;
  assign n32310 = ~n6056 & n32309;
  assign n32311 = ~n7073 & n32310;
  assign n32312 = ~n8179 & n32311;
  assign n32313 = ~n9344 & n32312;
  assign n32314 = ~n13517 & n32313;
  assign n32315 = ~n13516 & n32314;
  assign n32316 = ~n10594 & n32315;
  assign n32317 = ~n12861 & n32316;
  assign n32318 = ~n12005 & n32317;
  assign n32319 = ~n13515 & n32318;
  assign n32320 = n13532 & n32319;
  assign n32321 = n13514 & n32320;
  assign n32322 = n13557 & n32321;
  assign n32323 = ~n32305 & ~n32322;
  assign n32324 = ~n32289 & n32323;
  assign n32325 = pi186 & ~n9717;
  assign n32326 = ~n9913 & n32325;
  assign n32327 = n9856 & n32326;
  assign n32328 = ~n9929 & n32327;
  assign n32329 = ~n13824 & n32328;
  assign n32330 = ~n13823 & n32329;
  assign n32331 = ~n11266 & n32330;
  assign n32332 = ~n12861 & n32331;
  assign n32333 = ~n11588 & n32332;
  assign n32334 = ~n12973 & n32333;
  assign n32335 = n13054 & n32334;
  assign n32336 = n13095 & n32335;
  assign n32337 = n13858 & n32336;
  assign n32338 = pi218 & ~n12671;
  assign n32339 = ~n12811 & n32338;
  assign n32340 = n13912 & n32339;
  assign n32341 = ~n12902 & n32340;
  assign n32342 = ~n13908 & n32341;
  assign n32343 = ~n12861 & n32342;
  assign n32344 = ~n12860 & n32343;
  assign n32345 = n12952 & n32344;
  assign n32346 = n13919 & n32345;
  assign n32347 = n14008 & n32346;
  assign n32348 = ~n32337 & ~n32347;
  assign n32349 = ~n12861 & n29864;
  assign n32350 = ~n12471 & n32349;
  assign n32351 = ~n12972 & n32350;
  assign n32352 = n14020 & n32351;
  assign n32353 = n13095 & n32352;
  assign n32354 = n14072 & n32353;
  assign n32355 = pi202 & ~n10909;
  assign n32356 = ~n11168 & n32355;
  assign n32357 = n11135 & n32356;
  assign n32358 = ~n11188 & n32357;
  assign n32359 = ~n14011 & n32358;
  assign n32360 = ~n14010 & n32359;
  assign n32361 = ~n12861 & n32360;
  assign n32362 = ~n12380 & n32361;
  assign n32363 = ~n12972 & n32362;
  assign n32364 = n14020 & n32363;
  assign n32365 = n13095 & n32364;
  assign n32366 = n14044 & n32365;
  assign n32367 = ~n32354 & ~n32366;
  assign n32368 = n32348 & n32367;
  assign n32369 = n13319 & n25413;
  assign n32370 = ~n3066 & n32369;
  assign n32371 = ~n3983 & n32370;
  assign n32372 = ~n4003 & n32371;
  assign n32373 = ~n4024 & n32372;
  assign n32374 = ~n4999 & n32373;
  assign n32375 = ~n5827 & n32374;
  assign n32376 = ~n6893 & n32375;
  assign n32377 = ~n7890 & n32376;
  assign n32378 = ~n9131 & n32377;
  assign n32379 = ~n13144 & n32378;
  assign n32380 = ~n13143 & n32379;
  assign n32381 = ~n10278 & n32380;
  assign n32382 = ~n13142 & n32381;
  assign n32383 = ~n11662 & n32382;
  assign n32384 = ~n13141 & n32383;
  assign n32385 = n13165 & n32384;
  assign n32386 = n13140 & n32385;
  assign n32387 = n13190 & n32386;
  assign n32388 = pi226 & ~n12946;
  assign n32389 = ~n12903 & n32388;
  assign n32390 = ~n12861 & n32389;
  assign n32391 = ~n12860 & n32390;
  assign n32392 = n12952 & n32391;
  assign n32393 = n12975 & n32392;
  assign n32394 = n13092 & n32393;
  assign n32395 = ~n32387 & ~n32394;
  assign n32396 = n13408 & n27507;
  assign n32397 = ~n3940 & n32396;
  assign n32398 = ~n4001 & n32397;
  assign n32399 = ~n5043 & n32398;
  assign n32400 = ~n5943 & n32399;
  assign n32401 = ~n6951 & n32400;
  assign n32402 = ~n8037 & n32401;
  assign n32403 = ~n9200 & n32402;
  assign n32404 = ~n13348 & n32403;
  assign n32405 = ~n13347 & n32404;
  assign n32406 = ~n10445 & n32405;
  assign n32407 = ~n12861 & n32406;
  assign n32408 = ~n11846 & n32407;
  assign n32409 = ~n13346 & n32408;
  assign n32410 = n13367 & n32409;
  assign n32411 = n13345 & n32410;
  assign n32412 = n13392 & n32411;
  assign n32413 = pi170 & ~n8574;
  assign n32414 = n11377 & n32413;
  assign n32415 = n9942 & n32414;
  assign n32416 = ~n8834 & n32415;
  assign n32417 = ~n10002 & n32416;
  assign n32418 = ~n13097 & n32417;
  assign n32419 = ~n13096 & n32418;
  assign n32420 = ~n11297 & n32419;
  assign n32421 = ~n12861 & n32420;
  assign n32422 = ~n12240 & n32421;
  assign n32423 = ~n12973 & n32422;
  assign n32424 = n13109 & n32423;
  assign n32425 = n13095 & n32424;
  assign n32426 = n13134 & n32425;
  assign n32427 = ~n32412 & ~n32426;
  assign n32428 = n32395 & n32427;
  assign n32429 = n32368 & n32428;
  assign n32430 = n32324 & n32429;
  assign po123 = ~n32274 | ~n32430;
  assign n32432 = ~n11343 & n30076;
  assign n32433 = ~n12861 & n32432;
  assign n32434 = ~n11551 & n32433;
  assign n32435 = ~n12973 & n32434;
  assign n32436 = n13095 & n32435;
  assign n32437 = n13885 & n32436;
  assign n32438 = n13905 & n32437;
  assign n32439 = ~n10705 & n30166;
  assign n32440 = ~n12861 & n32439;
  assign n32441 = ~n12121 & n32440;
  assign n32442 = ~n13717 & n32441;
  assign n32443 = n13723 & n32442;
  assign n32444 = n13095 & n32443;
  assign n32445 = n13716 & n32444;
  assign n32446 = ~n32438 & ~n32445;
  assign n32447 = ~n11318 & n30159;
  assign n32448 = ~n12861 & n32447;
  assign n32449 = ~n12181 & n32448;
  assign n32450 = ~n13052 & n32449;
  assign n32451 = n13095 & n32450;
  assign n32452 = n13758 & n32451;
  assign n32453 = n13751 & n32452;
  assign n32454 = ~n10787 & n30137;
  assign n32455 = ~n12861 & n32454;
  assign n32456 = ~n11611 & n32455;
  assign n32457 = ~n12973 & n32456;
  assign n32458 = n13802 & n32457;
  assign n32459 = n13095 & n32458;
  assign n32460 = n13819 & n32459;
  assign n32461 = ~n32453 & ~n32460;
  assign n32462 = n32446 & n32461;
  assign n32463 = pi059 & ~n1679;
  assign n32464 = n1741 & n32463;
  assign n32465 = n13259 & n32464;
  assign n32466 = ~n2242 & n32465;
  assign n32467 = ~n3095 & n32466;
  assign n32468 = ~n3997 & n32467;
  assign n32469 = ~n4003 & n32468;
  assign n32470 = ~n4837 & n32469;
  assign n32471 = ~n5822 & n32470;
  assign n32472 = ~n6820 & n32471;
  assign n32473 = ~n7785 & n32472;
  assign n32474 = ~n9027 & n32473;
  assign n32475 = ~n10245 & n32474;
  assign n32476 = ~n13258 & n32475;
  assign n32477 = ~n13257 & n32476;
  assign n32478 = ~n11536 & n32477;
  assign n32479 = ~n13256 & n32478;
  assign n32480 = ~n13036 & n32479;
  assign n32481 = ~n13255 & n32480;
  assign n32482 = n13281 & n32481;
  assign n32483 = n13254 & n32482;
  assign n32484 = n13306 & n32483;
  assign n32485 = ~n11860 & n29877;
  assign n32486 = ~n12861 & n32485;
  assign n32487 = ~n13399 & n32486;
  assign n32488 = n13406 & n32487;
  assign n32489 = ~n13312 & n29881;
  assign n32490 = ~n13310 & n32489;
  assign n32491 = n13317 & n32490;
  assign n32492 = pi243 & ~n501;
  assign n32493 = n14188 & n32492;
  assign n32494 = n31189 & n32493;
  assign n32495 = n31196 & n32494;
  assign n32496 = ~n1172 & n32495;
  assign n32497 = ~n996 & n32496;
  assign n32498 = ~n2306 & n32497;
  assign n32499 = n3819 & n32498;
  assign n32500 = n3821 & n32499;
  assign n32501 = n14186 & n32500;
  assign n32502 = n14229 & n32501;
  assign n32503 = n14184 & n32502;
  assign n32504 = n14180 & n32503;
  assign n32505 = ~n7236 & n32504;
  assign n32506 = ~n6137 & n32505;
  assign n32507 = n6193 & n32506;
  assign n32508 = n6134 & n32507;
  assign n32509 = ~n8867 & n32508;
  assign n32510 = ~n7235 & n32509;
  assign n32511 = n7296 & n32510;
  assign n32512 = n7231 & n32511;
  assign n32513 = ~n10027 & n32512;
  assign n32514 = ~n8866 & n32513;
  assign n32515 = n8898 & n32514;
  assign n32516 = n8863 & n32515;
  assign n32517 = pi235 & ~n501;
  assign n32518 = n14255 & n32517;
  assign n32519 = n14253 & n32518;
  assign n32520 = n31154 & n32519;
  assign n32521 = n31162 & n32520;
  assign n32522 = ~n1172 & n32521;
  assign n32523 = ~n996 & n32522;
  assign n32524 = ~n2306 & n32523;
  assign n32525 = n3819 & n32524;
  assign n32526 = n14139 & n32525;
  assign n32527 = n12583 & n32526;
  assign n32528 = n14252 & n32527;
  assign n32529 = n14242 & n32528;
  assign n32530 = n14431 & n32529;
  assign n32531 = ~n7236 & n32530;
  assign n32532 = ~n6137 & n32531;
  assign n32533 = n6193 & n32532;
  assign n32534 = n6134 & n32533;
  assign n32535 = ~n8867 & n32534;
  assign n32536 = ~n7235 & n32535;
  assign n32537 = n7296 & n32536;
  assign n32538 = n7231 & n32537;
  assign n32539 = ~n10027 & n32538;
  assign n32540 = ~n8866 & n32539;
  assign n32541 = n8898 & n32540;
  assign n32542 = n8863 & n32541;
  assign n32543 = ~n32516 & ~n32542;
  assign n32544 = ~n10788 & ~n32543;
  assign n32545 = ~n10026 & n32544;
  assign n32546 = n10072 & n32545;
  assign n32547 = n10021 & n32546;
  assign n32548 = ~n32491 & ~n32547;
  assign n32549 = ~n32488 & n32548;
  assign n32550 = ~n11959 & n29945;
  assign n32551 = ~n12861 & n32550;
  assign n32552 = ~n12950 & n32551;
  assign n32553 = n13491 & n32552;
  assign n32554 = n13486 & n32553;
  assign n32555 = ~n12041 & n29950;
  assign n32556 = ~n12861 & n32555;
  assign n32557 = n13094 & n32556;
  assign n32558 = n13577 & n32557;
  assign n32559 = n13572 & n32558;
  assign n32560 = ~n32554 & ~n32559;
  assign n32561 = n32549 & n32560;
  assign n32562 = ~n32484 & n32561;
  assign n32563 = n13731 & n25575;
  assign n32564 = ~n7869 & n32563;
  assign n32565 = ~n8346 & n32564;
  assign n32566 = ~n9485 & n32565;
  assign n32567 = ~n13653 & n32566;
  assign n32568 = ~n13652 & n32567;
  assign n32569 = ~n10741 & n32568;
  assign n32570 = ~n12861 & n32569;
  assign n32571 = ~n12158 & n32570;
  assign n32572 = ~n13052 & n32571;
  assign n32573 = n13667 & n32572;
  assign n32574 = n13095 & n32573;
  assign n32575 = n13692 & n32574;
  assign n32576 = pi227 & ~n12946;
  assign n32577 = ~n12903 & n32576;
  assign n32578 = ~n12861 & n32577;
  assign n32579 = ~n12860 & n32578;
  assign n32580 = n12952 & n32579;
  assign n32581 = n12975 & n32580;
  assign n32582 = n13092 & n32581;
  assign n32583 = ~n32575 & ~n32582;
  assign n32584 = n32562 & n32583;
  assign n32585 = n32462 & n32584;
  assign n32586 = pi123 & ~n5627;
  assign n32587 = n5687 & n32586;
  assign n32588 = n13580 & n32587;
  assign n32589 = ~n5808 & n32588;
  assign n32590 = ~n6056 & n32589;
  assign n32591 = ~n7073 & n32590;
  assign n32592 = ~n8179 & n32591;
  assign n32593 = ~n9344 & n32592;
  assign n32594 = ~n13517 & n32593;
  assign n32595 = ~n13516 & n32594;
  assign n32596 = ~n10594 & n32595;
  assign n32597 = ~n12861 & n32596;
  assign n32598 = ~n12005 & n32597;
  assign n32599 = ~n13515 & n32598;
  assign n32600 = n13532 & n32599;
  assign n32601 = n13514 & n32600;
  assign n32602 = n13557 & n32601;
  assign n32603 = n13408 & n27771;
  assign n32604 = ~n3940 & n32603;
  assign n32605 = ~n4001 & n32604;
  assign n32606 = ~n5043 & n32605;
  assign n32607 = ~n5943 & n32606;
  assign n32608 = ~n6951 & n32607;
  assign n32609 = ~n8037 & n32608;
  assign n32610 = ~n9200 & n32609;
  assign n32611 = ~n13348 & n32610;
  assign n32612 = ~n13347 & n32611;
  assign n32613 = ~n10445 & n32612;
  assign n32614 = ~n12861 & n32613;
  assign n32615 = ~n11846 & n32614;
  assign n32616 = ~n13346 & n32615;
  assign n32617 = n13367 & n32616;
  assign n32618 = n13345 & n32617;
  assign n32619 = n13392 & n32618;
  assign n32620 = n13494 & n27804;
  assign n32621 = ~n4817 & n32620;
  assign n32622 = ~n4902 & n32621;
  assign n32623 = ~n6001 & n32622;
  assign n32624 = ~n7014 & n32623;
  assign n32625 = ~n8114 & n32624;
  assign n32626 = ~n9276 & n32625;
  assign n32627 = ~n13438 & n32626;
  assign n32628 = ~n13437 & n32627;
  assign n32629 = ~n10523 & n32628;
  assign n32630 = ~n12861 & n32629;
  assign n32631 = ~n11928 & n32630;
  assign n32632 = ~n13436 & n32631;
  assign n32633 = n13453 & n32632;
  assign n32634 = n13435 & n32633;
  assign n32635 = n13478 & n32634;
  assign n32636 = ~n32619 & ~n32635;
  assign n32637 = ~n32602 & n32636;
  assign n32638 = ~n12861 & n30085;
  assign n32639 = ~n12471 & n32638;
  assign n32640 = ~n12972 & n32639;
  assign n32641 = n14020 & n32640;
  assign n32642 = n13095 & n32641;
  assign n32643 = n14072 & n32642;
  assign n32644 = n13319 & n25670;
  assign n32645 = ~n3066 & n32644;
  assign n32646 = ~n3983 & n32645;
  assign n32647 = ~n4003 & n32646;
  assign n32648 = ~n4024 & n32647;
  assign n32649 = ~n4999 & n32648;
  assign n32650 = ~n5827 & n32649;
  assign n32651 = ~n6893 & n32650;
  assign n32652 = ~n7890 & n32651;
  assign n32653 = ~n9131 & n32652;
  assign n32654 = ~n13144 & n32653;
  assign n32655 = ~n13143 & n32654;
  assign n32656 = ~n10278 & n32655;
  assign n32657 = ~n13142 & n32656;
  assign n32658 = ~n11662 & n32657;
  assign n32659 = ~n13141 & n32658;
  assign n32660 = n13165 & n32659;
  assign n32661 = n13140 & n32660;
  assign n32662 = n13190 & n32661;
  assign n32663 = ~n32643 & ~n32662;
  assign n32664 = n13202 & n27732;
  assign n32665 = ~n1372 & n32664;
  assign n32666 = ~n2243 & n32665;
  assign n32667 = ~n3104 & n32666;
  assign n32668 = ~n3971 & n32667;
  assign n32669 = ~n4003 & n32668;
  assign n32670 = ~n4872 & n32669;
  assign n32671 = ~n5801 & n32670;
  assign n32672 = ~n6739 & n32671;
  assign n32673 = ~n7807 & n32672;
  assign n32674 = ~n8989 & n32673;
  assign n32675 = ~n10273 & n32674;
  assign n32676 = ~n13200 & n32675;
  assign n32677 = ~n13199 & n32676;
  assign n32678 = ~n11499 & n32677;
  assign n32679 = ~n13198 & n32678;
  assign n32680 = ~n13076 & n32679;
  assign n32681 = ~n13197 & n32680;
  assign n32682 = n13223 & n32681;
  assign n32683 = n13196 & n32682;
  assign n32684 = n13248 & n32683;
  assign n32685 = n7175 & n27789;
  assign n32686 = n13694 & n32685;
  assign n32687 = ~n6784 & n32686;
  assign n32688 = ~n7158 & n32687;
  assign n32689 = ~n8250 & n32688;
  assign n32690 = ~n9414 & n32689;
  assign n32691 = ~n13602 & n32690;
  assign n32692 = ~n13601 & n32691;
  assign n32693 = ~n10667 & n32692;
  assign n32694 = ~n12861 & n32693;
  assign n32695 = ~n12083 & n32694;
  assign n32696 = ~n13600 & n32695;
  assign n32697 = n13618 & n32696;
  assign n32698 = n13095 & n32697;
  assign n32699 = n13643 & n32698;
  assign n32700 = ~n32684 & ~n32699;
  assign n32701 = n32663 & n32700;
  assign n32702 = pi203 & ~n10909;
  assign n32703 = ~n11168 & n32702;
  assign n32704 = n11135 & n32703;
  assign n32705 = ~n11188 & n32704;
  assign n32706 = ~n14011 & n32705;
  assign n32707 = ~n14010 & n32706;
  assign n32708 = ~n12861 & n32707;
  assign n32709 = ~n12380 & n32708;
  assign n32710 = ~n12972 & n32709;
  assign n32711 = n14020 & n32710;
  assign n32712 = n13095 & n32711;
  assign n32713 = n14044 & n32712;
  assign n32714 = pi219 & ~n12671;
  assign n32715 = ~n12811 & n32714;
  assign n32716 = n13912 & n32715;
  assign n32717 = ~n12902 & n32716;
  assign n32718 = ~n13908 & n32717;
  assign n32719 = ~n12861 & n32718;
  assign n32720 = ~n12860 & n32719;
  assign n32721 = n12952 & n32720;
  assign n32722 = n13919 & n32721;
  assign n32723 = n14008 & n32722;
  assign n32724 = ~n32713 & ~n32723;
  assign n32725 = pi171 & ~n8574;
  assign n32726 = n11377 & n32725;
  assign n32727 = n9942 & n32726;
  assign n32728 = ~n8834 & n32727;
  assign n32729 = ~n10002 & n32728;
  assign n32730 = ~n13097 & n32729;
  assign n32731 = ~n13096 & n32730;
  assign n32732 = ~n11297 & n32731;
  assign n32733 = ~n12861 & n32732;
  assign n32734 = ~n12240 & n32733;
  assign n32735 = ~n12973 & n32734;
  assign n32736 = n13109 & n32735;
  assign n32737 = n13095 & n32736;
  assign n32738 = n13134 & n32737;
  assign n32739 = pi187 & ~n9717;
  assign n32740 = ~n9913 & n32739;
  assign n32741 = n9856 & n32740;
  assign n32742 = ~n9929 & n32741;
  assign n32743 = ~n13824 & n32742;
  assign n32744 = ~n13823 & n32743;
  assign n32745 = ~n11266 & n32744;
  assign n32746 = ~n12861 & n32745;
  assign n32747 = ~n11588 & n32746;
  assign n32748 = ~n12973 & n32747;
  assign n32749 = n13054 & n32748;
  assign n32750 = n13095 & n32749;
  assign n32751 = n13858 & n32750;
  assign n32752 = ~n32738 & ~n32751;
  assign n32753 = n32724 & n32752;
  assign n32754 = n32701 & n32753;
  assign n32755 = n32637 & n32754;
  assign po124 = ~n32585 | ~n32755;
  assign n32757 = ~n10705 & n30467;
  assign n32758 = ~n12861 & n32757;
  assign n32759 = ~n12121 & n32758;
  assign n32760 = ~n13717 & n32759;
  assign n32761 = n13723 & n32760;
  assign n32762 = n13095 & n32761;
  assign n32763 = n13716 & n32762;
  assign n32764 = ~n11318 & n30460;
  assign n32765 = ~n12861 & n32764;
  assign n32766 = ~n12181 & n32765;
  assign n32767 = ~n13052 & n32766;
  assign n32768 = n13095 & n32767;
  assign n32769 = n13758 & n32768;
  assign n32770 = n13751 & n32769;
  assign n32771 = ~n32763 & ~n32770;
  assign n32772 = ~n10787 & n30438;
  assign n32773 = ~n12861 & n32772;
  assign n32774 = ~n11611 & n32773;
  assign n32775 = ~n12973 & n32774;
  assign n32776 = n13802 & n32775;
  assign n32777 = n13095 & n32776;
  assign n32778 = n13819 & n32777;
  assign n32779 = ~n11343 & n30377;
  assign n32780 = ~n12861 & n32779;
  assign n32781 = ~n11551 & n32780;
  assign n32782 = ~n12973 & n32781;
  assign n32783 = n13095 & n32782;
  assign n32784 = n13885 & n32783;
  assign n32785 = n13905 & n32784;
  assign n32786 = ~n32778 & ~n32785;
  assign n32787 = n32771 & n32786;
  assign n32788 = n13731 & n25808;
  assign n32789 = ~n7869 & n32788;
  assign n32790 = ~n8346 & n32789;
  assign n32791 = ~n9485 & n32790;
  assign n32792 = ~n13653 & n32791;
  assign n32793 = ~n13652 & n32792;
  assign n32794 = ~n10741 & n32793;
  assign n32795 = ~n12861 & n32794;
  assign n32796 = ~n12158 & n32795;
  assign n32797 = ~n13052 & n32796;
  assign n32798 = n13667 & n32797;
  assign n32799 = n13095 & n32798;
  assign n32800 = n13692 & n32799;
  assign n32801 = ~n11860 & n30178;
  assign n32802 = ~n12861 & n32801;
  assign n32803 = ~n13399 & n32802;
  assign n32804 = n13406 & n32803;
  assign n32805 = ~n13312 & n30182;
  assign n32806 = ~n13310 & n32805;
  assign n32807 = n13317 & n32806;
  assign n32808 = pi244 & ~n501;
  assign n32809 = n14188 & n32808;
  assign n32810 = n31189 & n32809;
  assign n32811 = n31196 & n32810;
  assign n32812 = ~n1172 & n32811;
  assign n32813 = ~n996 & n32812;
  assign n32814 = ~n2306 & n32813;
  assign n32815 = n3819 & n32814;
  assign n32816 = n3821 & n32815;
  assign n32817 = n14186 & n32816;
  assign n32818 = n14229 & n32817;
  assign n32819 = n14184 & n32818;
  assign n32820 = n14180 & n32819;
  assign n32821 = ~n7236 & n32820;
  assign n32822 = ~n6137 & n32821;
  assign n32823 = n6193 & n32822;
  assign n32824 = n6134 & n32823;
  assign n32825 = ~n8867 & n32824;
  assign n32826 = ~n7235 & n32825;
  assign n32827 = n7296 & n32826;
  assign n32828 = n7231 & n32827;
  assign n32829 = ~n10027 & n32828;
  assign n32830 = ~n8866 & n32829;
  assign n32831 = n8898 & n32830;
  assign n32832 = n8863 & n32831;
  assign n32833 = pi236 & ~n501;
  assign n32834 = n14255 & n32833;
  assign n32835 = n14253 & n32834;
  assign n32836 = n31154 & n32835;
  assign n32837 = n31162 & n32836;
  assign n32838 = ~n1172 & n32837;
  assign n32839 = ~n996 & n32838;
  assign n32840 = ~n2306 & n32839;
  assign n32841 = n3819 & n32840;
  assign n32842 = n14139 & n32841;
  assign n32843 = n12583 & n32842;
  assign n32844 = n14252 & n32843;
  assign n32845 = n14242 & n32844;
  assign n32846 = n14431 & n32845;
  assign n32847 = ~n7236 & n32846;
  assign n32848 = ~n6137 & n32847;
  assign n32849 = n6193 & n32848;
  assign n32850 = n6134 & n32849;
  assign n32851 = ~n8867 & n32850;
  assign n32852 = ~n7235 & n32851;
  assign n32853 = n7296 & n32852;
  assign n32854 = n7231 & n32853;
  assign n32855 = ~n10027 & n32854;
  assign n32856 = ~n8866 & n32855;
  assign n32857 = n8898 & n32856;
  assign n32858 = n8863 & n32857;
  assign n32859 = ~n32832 & ~n32858;
  assign n32860 = ~n10788 & ~n32859;
  assign n32861 = ~n10026 & n32860;
  assign n32862 = n10072 & n32861;
  assign n32863 = n10021 & n32862;
  assign n32864 = ~n32807 & ~n32863;
  assign n32865 = ~n32804 & n32864;
  assign n32866 = ~n11959 & n30246;
  assign n32867 = ~n12861 & n32866;
  assign n32868 = ~n12950 & n32867;
  assign n32869 = n13491 & n32868;
  assign n32870 = n13486 & n32869;
  assign n32871 = ~n12041 & n30251;
  assign n32872 = ~n12861 & n32871;
  assign n32873 = n13094 & n32872;
  assign n32874 = n13577 & n32873;
  assign n32875 = n13572 & n32874;
  assign n32876 = ~n32870 & ~n32875;
  assign n32877 = n32865 & n32876;
  assign n32878 = ~n32800 & n32877;
  assign n32879 = pi060 & ~n1679;
  assign n32880 = n1741 & n32879;
  assign n32881 = n13259 & n32880;
  assign n32882 = ~n2242 & n32881;
  assign n32883 = ~n3095 & n32882;
  assign n32884 = ~n3997 & n32883;
  assign n32885 = ~n4003 & n32884;
  assign n32886 = ~n4837 & n32885;
  assign n32887 = ~n5822 & n32886;
  assign n32888 = ~n6820 & n32887;
  assign n32889 = ~n7785 & n32888;
  assign n32890 = ~n9027 & n32889;
  assign n32891 = ~n10245 & n32890;
  assign n32892 = ~n13258 & n32891;
  assign n32893 = ~n13257 & n32892;
  assign n32894 = ~n11536 & n32893;
  assign n32895 = ~n13256 & n32894;
  assign n32896 = ~n13036 & n32895;
  assign n32897 = ~n13255 & n32896;
  assign n32898 = n13281 & n32897;
  assign n32899 = n13254 & n32898;
  assign n32900 = n13306 & n32899;
  assign n32901 = n13202 & n27998;
  assign n32902 = ~n1372 & n32901;
  assign n32903 = ~n2243 & n32902;
  assign n32904 = ~n3104 & n32903;
  assign n32905 = ~n3971 & n32904;
  assign n32906 = ~n4003 & n32905;
  assign n32907 = ~n4872 & n32906;
  assign n32908 = ~n5801 & n32907;
  assign n32909 = ~n6739 & n32908;
  assign n32910 = ~n7807 & n32909;
  assign n32911 = ~n8989 & n32910;
  assign n32912 = ~n10273 & n32911;
  assign n32913 = ~n13200 & n32912;
  assign n32914 = ~n13199 & n32913;
  assign n32915 = ~n11499 & n32914;
  assign n32916 = ~n13198 & n32915;
  assign n32917 = ~n13076 & n32916;
  assign n32918 = ~n13197 & n32917;
  assign n32919 = n13223 & n32918;
  assign n32920 = n13196 & n32919;
  assign n32921 = n13248 & n32920;
  assign n32922 = ~n32900 & ~n32921;
  assign n32923 = n32878 & n32922;
  assign n32924 = n32787 & n32923;
  assign n32925 = pi228 & ~n12946;
  assign n32926 = ~n12903 & n32925;
  assign n32927 = ~n12861 & n32926;
  assign n32928 = ~n12860 & n32927;
  assign n32929 = n12952 & n32928;
  assign n32930 = n12975 & n32929;
  assign n32931 = n13092 & n32930;
  assign n32932 = n7175 & n28055;
  assign n32933 = n13694 & n32932;
  assign n32934 = ~n6784 & n32933;
  assign n32935 = ~n7158 & n32934;
  assign n32936 = ~n8250 & n32935;
  assign n32937 = ~n9414 & n32936;
  assign n32938 = ~n13602 & n32937;
  assign n32939 = ~n13601 & n32938;
  assign n32940 = ~n10667 & n32939;
  assign n32941 = ~n12861 & n32940;
  assign n32942 = ~n12083 & n32941;
  assign n32943 = ~n13600 & n32942;
  assign n32944 = n13618 & n32943;
  assign n32945 = n13095 & n32944;
  assign n32946 = n13643 & n32945;
  assign n32947 = pi204 & ~n10909;
  assign n32948 = ~n11168 & n32947;
  assign n32949 = n11135 & n32948;
  assign n32950 = ~n11188 & n32949;
  assign n32951 = ~n14011 & n32950;
  assign n32952 = ~n14010 & n32951;
  assign n32953 = ~n12861 & n32952;
  assign n32954 = ~n12380 & n32953;
  assign n32955 = ~n12972 & n32954;
  assign n32956 = n14020 & n32955;
  assign n32957 = n13095 & n32956;
  assign n32958 = n14044 & n32957;
  assign n32959 = ~n32946 & ~n32958;
  assign n32960 = ~n32931 & n32959;
  assign n32961 = pi188 & ~n9717;
  assign n32962 = ~n9913 & n32961;
  assign n32963 = n9856 & n32962;
  assign n32964 = ~n9929 & n32963;
  assign n32965 = ~n13824 & n32964;
  assign n32966 = ~n13823 & n32965;
  assign n32967 = ~n11266 & n32966;
  assign n32968 = ~n12861 & n32967;
  assign n32969 = ~n11588 & n32968;
  assign n32970 = ~n12973 & n32969;
  assign n32971 = n13054 & n32970;
  assign n32972 = n13095 & n32971;
  assign n32973 = n13858 & n32972;
  assign n32974 = pi172 & ~n8574;
  assign n32975 = n11377 & n32974;
  assign n32976 = n9942 & n32975;
  assign n32977 = ~n8834 & n32976;
  assign n32978 = ~n10002 & n32977;
  assign n32979 = ~n13097 & n32978;
  assign n32980 = ~n13096 & n32979;
  assign n32981 = ~n11297 & n32980;
  assign n32982 = ~n12861 & n32981;
  assign n32983 = ~n12240 & n32982;
  assign n32984 = ~n12973 & n32983;
  assign n32985 = n13109 & n32984;
  assign n32986 = n13095 & n32985;
  assign n32987 = n13134 & n32986;
  assign n32988 = ~n32973 & ~n32987;
  assign n32989 = pi124 & ~n5627;
  assign n32990 = n5687 & n32989;
  assign n32991 = n13580 & n32990;
  assign n32992 = ~n5808 & n32991;
  assign n32993 = ~n6056 & n32992;
  assign n32994 = ~n7073 & n32993;
  assign n32995 = ~n8179 & n32994;
  assign n32996 = ~n9344 & n32995;
  assign n32997 = ~n13517 & n32996;
  assign n32998 = ~n13516 & n32997;
  assign n32999 = ~n10594 & n32998;
  assign n33000 = ~n12861 & n32999;
  assign n33001 = ~n12005 & n33000;
  assign n33002 = ~n13515 & n33001;
  assign n33003 = n13532 & n33002;
  assign n33004 = n13514 & n33003;
  assign n33005 = n13557 & n33004;
  assign n33006 = pi220 & ~n12671;
  assign n33007 = ~n12811 & n33006;
  assign n33008 = n13912 & n33007;
  assign n33009 = ~n12902 & n33008;
  assign n33010 = ~n13908 & n33009;
  assign n33011 = ~n12861 & n33010;
  assign n33012 = ~n12860 & n33011;
  assign n33013 = n12952 & n33012;
  assign n33014 = n13919 & n33013;
  assign n33015 = n14008 & n33014;
  assign n33016 = ~n33005 & ~n33015;
  assign n33017 = n32988 & n33016;
  assign n33018 = n13408 & n28037;
  assign n33019 = ~n3940 & n33018;
  assign n33020 = ~n4001 & n33019;
  assign n33021 = ~n5043 & n33020;
  assign n33022 = ~n5943 & n33021;
  assign n33023 = ~n6951 & n33022;
  assign n33024 = ~n8037 & n33023;
  assign n33025 = ~n9200 & n33024;
  assign n33026 = ~n13348 & n33025;
  assign n33027 = ~n13347 & n33026;
  assign n33028 = ~n10445 & n33027;
  assign n33029 = ~n12861 & n33028;
  assign n33030 = ~n11846 & n33029;
  assign n33031 = ~n13346 & n33030;
  assign n33032 = n13367 & n33031;
  assign n33033 = n13345 & n33032;
  assign n33034 = n13392 & n33033;
  assign n33035 = n13319 & n25903;
  assign n33036 = ~n3066 & n33035;
  assign n33037 = ~n3983 & n33036;
  assign n33038 = ~n4003 & n33037;
  assign n33039 = ~n4024 & n33038;
  assign n33040 = ~n4999 & n33039;
  assign n33041 = ~n5827 & n33040;
  assign n33042 = ~n6893 & n33041;
  assign n33043 = ~n7890 & n33042;
  assign n33044 = ~n9131 & n33043;
  assign n33045 = ~n13144 & n33044;
  assign n33046 = ~n13143 & n33045;
  assign n33047 = ~n10278 & n33046;
  assign n33048 = ~n13142 & n33047;
  assign n33049 = ~n11662 & n33048;
  assign n33050 = ~n13141 & n33049;
  assign n33051 = n13165 & n33050;
  assign n33052 = n13140 & n33051;
  assign n33053 = n13190 & n33052;
  assign n33054 = ~n33034 & ~n33053;
  assign n33055 = ~n12861 & n30386;
  assign n33056 = ~n12471 & n33055;
  assign n33057 = ~n12972 & n33056;
  assign n33058 = n14020 & n33057;
  assign n33059 = n13095 & n33058;
  assign n33060 = n14072 & n33059;
  assign n33061 = n13494 & n28070;
  assign n33062 = ~n4817 & n33061;
  assign n33063 = ~n4902 & n33062;
  assign n33064 = ~n6001 & n33063;
  assign n33065 = ~n7014 & n33064;
  assign n33066 = ~n8114 & n33065;
  assign n33067 = ~n9276 & n33066;
  assign n33068 = ~n13438 & n33067;
  assign n33069 = ~n13437 & n33068;
  assign n33070 = ~n10523 & n33069;
  assign n33071 = ~n12861 & n33070;
  assign n33072 = ~n11928 & n33071;
  assign n33073 = ~n13436 & n33072;
  assign n33074 = n13453 & n33073;
  assign n33075 = n13435 & n33074;
  assign n33076 = n13478 & n33075;
  assign n33077 = ~n33060 & ~n33076;
  assign n33078 = n33054 & n33077;
  assign n33079 = n33017 & n33078;
  assign n33080 = n32960 & n33079;
  assign po125 = ~n32924 | ~n33080;
  assign n33082 = ~n10705 & n30768;
  assign n33083 = ~n12861 & n33082;
  assign n33084 = ~n12121 & n33083;
  assign n33085 = ~n13717 & n33084;
  assign n33086 = n13723 & n33085;
  assign n33087 = n13095 & n33086;
  assign n33088 = n13716 & n33087;
  assign n33089 = ~n11318 & n30761;
  assign n33090 = ~n12861 & n33089;
  assign n33091 = ~n12181 & n33090;
  assign n33092 = ~n13052 & n33091;
  assign n33093 = n13095 & n33092;
  assign n33094 = n13758 & n33093;
  assign n33095 = n13751 & n33094;
  assign n33096 = ~n33088 & ~n33095;
  assign n33097 = ~n10787 & n30739;
  assign n33098 = ~n12861 & n33097;
  assign n33099 = ~n11611 & n33098;
  assign n33100 = ~n12973 & n33099;
  assign n33101 = n13802 & n33100;
  assign n33102 = n13095 & n33101;
  assign n33103 = n13819 & n33102;
  assign n33104 = ~n11343 & n30678;
  assign n33105 = ~n12861 & n33104;
  assign n33106 = ~n11551 & n33105;
  assign n33107 = ~n12973 & n33106;
  assign n33108 = n13095 & n33107;
  assign n33109 = n13885 & n33108;
  assign n33110 = n13905 & n33109;
  assign n33111 = ~n33103 & ~n33110;
  assign n33112 = n33096 & n33111;
  assign n33113 = n13731 & n26041;
  assign n33114 = ~n7869 & n33113;
  assign n33115 = ~n8346 & n33114;
  assign n33116 = ~n9485 & n33115;
  assign n33117 = ~n13653 & n33116;
  assign n33118 = ~n13652 & n33117;
  assign n33119 = ~n10741 & n33118;
  assign n33120 = ~n12861 & n33119;
  assign n33121 = ~n12158 & n33120;
  assign n33122 = ~n13052 & n33121;
  assign n33123 = n13667 & n33122;
  assign n33124 = n13095 & n33123;
  assign n33125 = n13692 & n33124;
  assign n33126 = ~n11860 & n30479;
  assign n33127 = ~n12861 & n33126;
  assign n33128 = ~n13399 & n33127;
  assign n33129 = n13406 & n33128;
  assign n33130 = ~n13312 & n30483;
  assign n33131 = ~n13310 & n33130;
  assign n33132 = n13317 & n33131;
  assign n33133 = pi237 & ~n501;
  assign n33134 = n14255 & n33133;
  assign n33135 = n14253 & n33134;
  assign n33136 = n31154 & n33135;
  assign n33137 = n31162 & n33136;
  assign n33138 = ~n1172 & n33137;
  assign n33139 = ~n996 & n33138;
  assign n33140 = ~n2306 & n33139;
  assign n33141 = n3819 & n33140;
  assign n33142 = n14139 & n33141;
  assign n33143 = n12583 & n33142;
  assign n33144 = n14252 & n33143;
  assign n33145 = n14242 & n33144;
  assign n33146 = n14431 & n33145;
  assign n33147 = ~n7236 & n33146;
  assign n33148 = ~n6137 & n33147;
  assign n33149 = n6193 & n33148;
  assign n33150 = n6134 & n33149;
  assign n33151 = ~n8867 & n33150;
  assign n33152 = ~n7235 & n33151;
  assign n33153 = n7296 & n33152;
  assign n33154 = n7231 & n33153;
  assign n33155 = ~n10027 & n33154;
  assign n33156 = ~n8866 & n33155;
  assign n33157 = n8898 & n33156;
  assign n33158 = n8863 & n33157;
  assign n33159 = pi245 & ~n501;
  assign n33160 = n14188 & n33159;
  assign n33161 = n31189 & n33160;
  assign n33162 = n31196 & n33161;
  assign n33163 = ~n1172 & n33162;
  assign n33164 = ~n996 & n33163;
  assign n33165 = ~n2306 & n33164;
  assign n33166 = n3819 & n33165;
  assign n33167 = n3821 & n33166;
  assign n33168 = n14186 & n33167;
  assign n33169 = n14229 & n33168;
  assign n33170 = n14184 & n33169;
  assign n33171 = n14180 & n33170;
  assign n33172 = ~n7236 & n33171;
  assign n33173 = ~n6137 & n33172;
  assign n33174 = n6193 & n33173;
  assign n33175 = n6134 & n33174;
  assign n33176 = ~n8867 & n33175;
  assign n33177 = ~n7235 & n33176;
  assign n33178 = n7296 & n33177;
  assign n33179 = n7231 & n33178;
  assign n33180 = ~n10027 & n33179;
  assign n33181 = ~n8866 & n33180;
  assign n33182 = n8898 & n33181;
  assign n33183 = n8863 & n33182;
  assign n33184 = ~n33158 & ~n33183;
  assign n33185 = ~n10788 & ~n33184;
  assign n33186 = ~n10026 & n33185;
  assign n33187 = n10072 & n33186;
  assign n33188 = n10021 & n33187;
  assign n33189 = ~n33132 & ~n33188;
  assign n33190 = ~n33129 & n33189;
  assign n33191 = ~n11959 & n30547;
  assign n33192 = ~n12861 & n33191;
  assign n33193 = ~n12950 & n33192;
  assign n33194 = n13491 & n33193;
  assign n33195 = n13486 & n33194;
  assign n33196 = ~n12041 & n30552;
  assign n33197 = ~n12861 & n33196;
  assign n33198 = n13094 & n33197;
  assign n33199 = n13577 & n33198;
  assign n33200 = n13572 & n33199;
  assign n33201 = ~n33195 & ~n33200;
  assign n33202 = n33190 & n33201;
  assign n33203 = ~n33125 & n33202;
  assign n33204 = pi061 & ~n1679;
  assign n33205 = n1741 & n33204;
  assign n33206 = n13259 & n33205;
  assign n33207 = ~n2242 & n33206;
  assign n33208 = ~n3095 & n33207;
  assign n33209 = ~n3997 & n33208;
  assign n33210 = ~n4003 & n33209;
  assign n33211 = ~n4837 & n33210;
  assign n33212 = ~n5822 & n33211;
  assign n33213 = ~n6820 & n33212;
  assign n33214 = ~n7785 & n33213;
  assign n33215 = ~n9027 & n33214;
  assign n33216 = ~n10245 & n33215;
  assign n33217 = ~n13258 & n33216;
  assign n33218 = ~n13257 & n33217;
  assign n33219 = ~n11536 & n33218;
  assign n33220 = ~n13256 & n33219;
  assign n33221 = ~n13036 & n33220;
  assign n33222 = ~n13255 & n33221;
  assign n33223 = n13281 & n33222;
  assign n33224 = n13254 & n33223;
  assign n33225 = n13306 & n33224;
  assign n33226 = n13202 & n28264;
  assign n33227 = ~n1372 & n33226;
  assign n33228 = ~n2243 & n33227;
  assign n33229 = ~n3104 & n33228;
  assign n33230 = ~n3971 & n33229;
  assign n33231 = ~n4003 & n33230;
  assign n33232 = ~n4872 & n33231;
  assign n33233 = ~n5801 & n33232;
  assign n33234 = ~n6739 & n33233;
  assign n33235 = ~n7807 & n33234;
  assign n33236 = ~n8989 & n33235;
  assign n33237 = ~n10273 & n33236;
  assign n33238 = ~n13200 & n33237;
  assign n33239 = ~n13199 & n33238;
  assign n33240 = ~n11499 & n33239;
  assign n33241 = ~n13198 & n33240;
  assign n33242 = ~n13076 & n33241;
  assign n33243 = ~n13197 & n33242;
  assign n33244 = n13223 & n33243;
  assign n33245 = n13196 & n33244;
  assign n33246 = n13248 & n33245;
  assign n33247 = ~n33225 & ~n33246;
  assign n33248 = n33203 & n33247;
  assign n33249 = n33112 & n33248;
  assign n33250 = pi229 & ~n12946;
  assign n33251 = ~n12903 & n33250;
  assign n33252 = ~n12861 & n33251;
  assign n33253 = ~n12860 & n33252;
  assign n33254 = n12952 & n33253;
  assign n33255 = n12975 & n33254;
  assign n33256 = n13092 & n33255;
  assign n33257 = n7175 & n28321;
  assign n33258 = n13694 & n33257;
  assign n33259 = ~n6784 & n33258;
  assign n33260 = ~n7158 & n33259;
  assign n33261 = ~n8250 & n33260;
  assign n33262 = ~n9414 & n33261;
  assign n33263 = ~n13602 & n33262;
  assign n33264 = ~n13601 & n33263;
  assign n33265 = ~n10667 & n33264;
  assign n33266 = ~n12861 & n33265;
  assign n33267 = ~n12083 & n33266;
  assign n33268 = ~n13600 & n33267;
  assign n33269 = n13618 & n33268;
  assign n33270 = n13095 & n33269;
  assign n33271 = n13643 & n33270;
  assign n33272 = pi205 & ~n10909;
  assign n33273 = ~n11168 & n33272;
  assign n33274 = n11135 & n33273;
  assign n33275 = ~n11188 & n33274;
  assign n33276 = ~n14011 & n33275;
  assign n33277 = ~n14010 & n33276;
  assign n33278 = ~n12861 & n33277;
  assign n33279 = ~n12380 & n33278;
  assign n33280 = ~n12972 & n33279;
  assign n33281 = n14020 & n33280;
  assign n33282 = n13095 & n33281;
  assign n33283 = n14044 & n33282;
  assign n33284 = ~n33271 & ~n33283;
  assign n33285 = ~n33256 & n33284;
  assign n33286 = pi189 & ~n9717;
  assign n33287 = ~n9913 & n33286;
  assign n33288 = n9856 & n33287;
  assign n33289 = ~n9929 & n33288;
  assign n33290 = ~n13824 & n33289;
  assign n33291 = ~n13823 & n33290;
  assign n33292 = ~n11266 & n33291;
  assign n33293 = ~n12861 & n33292;
  assign n33294 = ~n11588 & n33293;
  assign n33295 = ~n12973 & n33294;
  assign n33296 = n13054 & n33295;
  assign n33297 = n13095 & n33296;
  assign n33298 = n13858 & n33297;
  assign n33299 = pi173 & ~n8574;
  assign n33300 = n11377 & n33299;
  assign n33301 = n9942 & n33300;
  assign n33302 = ~n8834 & n33301;
  assign n33303 = ~n10002 & n33302;
  assign n33304 = ~n13097 & n33303;
  assign n33305 = ~n13096 & n33304;
  assign n33306 = ~n11297 & n33305;
  assign n33307 = ~n12861 & n33306;
  assign n33308 = ~n12240 & n33307;
  assign n33309 = ~n12973 & n33308;
  assign n33310 = n13109 & n33309;
  assign n33311 = n13095 & n33310;
  assign n33312 = n13134 & n33311;
  assign n33313 = ~n33298 & ~n33312;
  assign n33314 = pi125 & ~n5627;
  assign n33315 = n5687 & n33314;
  assign n33316 = n13580 & n33315;
  assign n33317 = ~n5808 & n33316;
  assign n33318 = ~n6056 & n33317;
  assign n33319 = ~n7073 & n33318;
  assign n33320 = ~n8179 & n33319;
  assign n33321 = ~n9344 & n33320;
  assign n33322 = ~n13517 & n33321;
  assign n33323 = ~n13516 & n33322;
  assign n33324 = ~n10594 & n33323;
  assign n33325 = ~n12861 & n33324;
  assign n33326 = ~n12005 & n33325;
  assign n33327 = ~n13515 & n33326;
  assign n33328 = n13532 & n33327;
  assign n33329 = n13514 & n33328;
  assign n33330 = n13557 & n33329;
  assign n33331 = pi221 & ~n12671;
  assign n33332 = ~n12811 & n33331;
  assign n33333 = n13912 & n33332;
  assign n33334 = ~n12902 & n33333;
  assign n33335 = ~n13908 & n33334;
  assign n33336 = ~n12861 & n33335;
  assign n33337 = ~n12860 & n33336;
  assign n33338 = n12952 & n33337;
  assign n33339 = n13919 & n33338;
  assign n33340 = n14008 & n33339;
  assign n33341 = ~n33330 & ~n33340;
  assign n33342 = n33313 & n33341;
  assign n33343 = n13408 & n28303;
  assign n33344 = ~n3940 & n33343;
  assign n33345 = ~n4001 & n33344;
  assign n33346 = ~n5043 & n33345;
  assign n33347 = ~n5943 & n33346;
  assign n33348 = ~n6951 & n33347;
  assign n33349 = ~n8037 & n33348;
  assign n33350 = ~n9200 & n33349;
  assign n33351 = ~n13348 & n33350;
  assign n33352 = ~n13347 & n33351;
  assign n33353 = ~n10445 & n33352;
  assign n33354 = ~n12861 & n33353;
  assign n33355 = ~n11846 & n33354;
  assign n33356 = ~n13346 & n33355;
  assign n33357 = n13367 & n33356;
  assign n33358 = n13345 & n33357;
  assign n33359 = n13392 & n33358;
  assign n33360 = n13319 & n26136;
  assign n33361 = ~n3066 & n33360;
  assign n33362 = ~n3983 & n33361;
  assign n33363 = ~n4003 & n33362;
  assign n33364 = ~n4024 & n33363;
  assign n33365 = ~n4999 & n33364;
  assign n33366 = ~n5827 & n33365;
  assign n33367 = ~n6893 & n33366;
  assign n33368 = ~n7890 & n33367;
  assign n33369 = ~n9131 & n33368;
  assign n33370 = ~n13144 & n33369;
  assign n33371 = ~n13143 & n33370;
  assign n33372 = ~n10278 & n33371;
  assign n33373 = ~n13142 & n33372;
  assign n33374 = ~n11662 & n33373;
  assign n33375 = ~n13141 & n33374;
  assign n33376 = n13165 & n33375;
  assign n33377 = n13140 & n33376;
  assign n33378 = n13190 & n33377;
  assign n33379 = ~n33359 & ~n33378;
  assign n33380 = ~n12861 & n30687;
  assign n33381 = ~n12471 & n33380;
  assign n33382 = ~n12972 & n33381;
  assign n33383 = n14020 & n33382;
  assign n33384 = n13095 & n33383;
  assign n33385 = n14072 & n33384;
  assign n33386 = n13494 & n28336;
  assign n33387 = ~n4817 & n33386;
  assign n33388 = ~n4902 & n33387;
  assign n33389 = ~n6001 & n33388;
  assign n33390 = ~n7014 & n33389;
  assign n33391 = ~n8114 & n33390;
  assign n33392 = ~n9276 & n33391;
  assign n33393 = ~n13438 & n33392;
  assign n33394 = ~n13437 & n33393;
  assign n33395 = ~n10523 & n33394;
  assign n33396 = ~n12861 & n33395;
  assign n33397 = ~n11928 & n33396;
  assign n33398 = ~n13436 & n33397;
  assign n33399 = n13453 & n33398;
  assign n33400 = n13435 & n33399;
  assign n33401 = n13478 & n33400;
  assign n33402 = ~n33385 & ~n33401;
  assign n33403 = n33379 & n33402;
  assign n33404 = n33342 & n33403;
  assign n33405 = n33285 & n33404;
  assign po126 = ~n33249 | ~n33405;
  assign n33407 = ~n10705 & n31069;
  assign n33408 = ~n12861 & n33407;
  assign n33409 = ~n12121 & n33408;
  assign n33410 = ~n13717 & n33409;
  assign n33411 = n13723 & n33410;
  assign n33412 = n13095 & n33411;
  assign n33413 = n13716 & n33412;
  assign n33414 = ~n11318 & n31062;
  assign n33415 = ~n12861 & n33414;
  assign n33416 = ~n12181 & n33415;
  assign n33417 = ~n13052 & n33416;
  assign n33418 = n13095 & n33417;
  assign n33419 = n13758 & n33418;
  assign n33420 = n13751 & n33419;
  assign n33421 = ~n33413 & ~n33420;
  assign n33422 = ~n10787 & n31040;
  assign n33423 = ~n12861 & n33422;
  assign n33424 = ~n11611 & n33423;
  assign n33425 = ~n12973 & n33424;
  assign n33426 = n13802 & n33425;
  assign n33427 = n13095 & n33426;
  assign n33428 = n13819 & n33427;
  assign n33429 = ~n11343 & n30979;
  assign n33430 = ~n12861 & n33429;
  assign n33431 = ~n11551 & n33430;
  assign n33432 = ~n12973 & n33431;
  assign n33433 = n13095 & n33432;
  assign n33434 = n13885 & n33433;
  assign n33435 = n13905 & n33434;
  assign n33436 = ~n33428 & ~n33435;
  assign n33437 = n33421 & n33436;
  assign n33438 = n13731 & n26274;
  assign n33439 = ~n7869 & n33438;
  assign n33440 = ~n8346 & n33439;
  assign n33441 = ~n9485 & n33440;
  assign n33442 = ~n13653 & n33441;
  assign n33443 = ~n13652 & n33442;
  assign n33444 = ~n10741 & n33443;
  assign n33445 = ~n12861 & n33444;
  assign n33446 = ~n12158 & n33445;
  assign n33447 = ~n13052 & n33446;
  assign n33448 = n13667 & n33447;
  assign n33449 = n13095 & n33448;
  assign n33450 = n13692 & n33449;
  assign n33451 = ~n11860 & n30780;
  assign n33452 = ~n12861 & n33451;
  assign n33453 = ~n13399 & n33452;
  assign n33454 = n13406 & n33453;
  assign n33455 = ~n13312 & n30784;
  assign n33456 = ~n13310 & n33455;
  assign n33457 = n13317 & n33456;
  assign n33458 = pi238 & ~n501;
  assign n33459 = n14255 & n33458;
  assign n33460 = n14253 & n33459;
  assign n33461 = n31154 & n33460;
  assign n33462 = n31162 & n33461;
  assign n33463 = ~n1172 & n33462;
  assign n33464 = ~n996 & n33463;
  assign n33465 = ~n2306 & n33464;
  assign n33466 = n3819 & n33465;
  assign n33467 = n14139 & n33466;
  assign n33468 = n12583 & n33467;
  assign n33469 = n14252 & n33468;
  assign n33470 = n14242 & n33469;
  assign n33471 = n14431 & n33470;
  assign n33472 = ~n7236 & n33471;
  assign n33473 = ~n6137 & n33472;
  assign n33474 = n6193 & n33473;
  assign n33475 = n6134 & n33474;
  assign n33476 = ~n8867 & n33475;
  assign n33477 = ~n7235 & n33476;
  assign n33478 = n7296 & n33477;
  assign n33479 = n7231 & n33478;
  assign n33480 = ~n10027 & n33479;
  assign n33481 = ~n8866 & n33480;
  assign n33482 = n8898 & n33481;
  assign n33483 = n8863 & n33482;
  assign n33484 = pi246 & ~n501;
  assign n33485 = n14188 & n33484;
  assign n33486 = n31189 & n33485;
  assign n33487 = n31196 & n33486;
  assign n33488 = ~n1172 & n33487;
  assign n33489 = ~n996 & n33488;
  assign n33490 = ~n2306 & n33489;
  assign n33491 = n3819 & n33490;
  assign n33492 = n3821 & n33491;
  assign n33493 = n14186 & n33492;
  assign n33494 = n14229 & n33493;
  assign n33495 = n14184 & n33494;
  assign n33496 = n14180 & n33495;
  assign n33497 = ~n7236 & n33496;
  assign n33498 = ~n6137 & n33497;
  assign n33499 = n6193 & n33498;
  assign n33500 = n6134 & n33499;
  assign n33501 = ~n8867 & n33500;
  assign n33502 = ~n7235 & n33501;
  assign n33503 = n7296 & n33502;
  assign n33504 = n7231 & n33503;
  assign n33505 = ~n10027 & n33504;
  assign n33506 = ~n8866 & n33505;
  assign n33507 = n8898 & n33506;
  assign n33508 = n8863 & n33507;
  assign n33509 = ~n33483 & ~n33508;
  assign n33510 = ~n10788 & ~n33509;
  assign n33511 = ~n10026 & n33510;
  assign n33512 = n10072 & n33511;
  assign n33513 = n10021 & n33512;
  assign n33514 = ~n33457 & ~n33513;
  assign n33515 = ~n33454 & n33514;
  assign n33516 = ~n11959 & n30848;
  assign n33517 = ~n12861 & n33516;
  assign n33518 = ~n12950 & n33517;
  assign n33519 = n13491 & n33518;
  assign n33520 = n13486 & n33519;
  assign n33521 = ~n12041 & n30853;
  assign n33522 = ~n12861 & n33521;
  assign n33523 = n13094 & n33522;
  assign n33524 = n13577 & n33523;
  assign n33525 = n13572 & n33524;
  assign n33526 = ~n33520 & ~n33525;
  assign n33527 = n33515 & n33526;
  assign n33528 = ~n33450 & n33527;
  assign n33529 = pi062 & ~n1679;
  assign n33530 = n1741 & n33529;
  assign n33531 = n13259 & n33530;
  assign n33532 = ~n2242 & n33531;
  assign n33533 = ~n3095 & n33532;
  assign n33534 = ~n3997 & n33533;
  assign n33535 = ~n4003 & n33534;
  assign n33536 = ~n4837 & n33535;
  assign n33537 = ~n5822 & n33536;
  assign n33538 = ~n6820 & n33537;
  assign n33539 = ~n7785 & n33538;
  assign n33540 = ~n9027 & n33539;
  assign n33541 = ~n10245 & n33540;
  assign n33542 = ~n13258 & n33541;
  assign n33543 = ~n13257 & n33542;
  assign n33544 = ~n11536 & n33543;
  assign n33545 = ~n13256 & n33544;
  assign n33546 = ~n13036 & n33545;
  assign n33547 = ~n13255 & n33546;
  assign n33548 = n13281 & n33547;
  assign n33549 = n13254 & n33548;
  assign n33550 = n13306 & n33549;
  assign n33551 = n13202 & n28530;
  assign n33552 = ~n1372 & n33551;
  assign n33553 = ~n2243 & n33552;
  assign n33554 = ~n3104 & n33553;
  assign n33555 = ~n3971 & n33554;
  assign n33556 = ~n4003 & n33555;
  assign n33557 = ~n4872 & n33556;
  assign n33558 = ~n5801 & n33557;
  assign n33559 = ~n6739 & n33558;
  assign n33560 = ~n7807 & n33559;
  assign n33561 = ~n8989 & n33560;
  assign n33562 = ~n10273 & n33561;
  assign n33563 = ~n13200 & n33562;
  assign n33564 = ~n13199 & n33563;
  assign n33565 = ~n11499 & n33564;
  assign n33566 = ~n13198 & n33565;
  assign n33567 = ~n13076 & n33566;
  assign n33568 = ~n13197 & n33567;
  assign n33569 = n13223 & n33568;
  assign n33570 = n13196 & n33569;
  assign n33571 = n13248 & n33570;
  assign n33572 = ~n33550 & ~n33571;
  assign n33573 = n33528 & n33572;
  assign n33574 = n33437 & n33573;
  assign n33575 = pi230 & ~n12946;
  assign n33576 = ~n12903 & n33575;
  assign n33577 = ~n12861 & n33576;
  assign n33578 = ~n12860 & n33577;
  assign n33579 = n12952 & n33578;
  assign n33580 = n12975 & n33579;
  assign n33581 = n13092 & n33580;
  assign n33582 = n7175 & n28587;
  assign n33583 = n13694 & n33582;
  assign n33584 = ~n6784 & n33583;
  assign n33585 = ~n7158 & n33584;
  assign n33586 = ~n8250 & n33585;
  assign n33587 = ~n9414 & n33586;
  assign n33588 = ~n13602 & n33587;
  assign n33589 = ~n13601 & n33588;
  assign n33590 = ~n10667 & n33589;
  assign n33591 = ~n12861 & n33590;
  assign n33592 = ~n12083 & n33591;
  assign n33593 = ~n13600 & n33592;
  assign n33594 = n13618 & n33593;
  assign n33595 = n13095 & n33594;
  assign n33596 = n13643 & n33595;
  assign n33597 = pi206 & ~n10909;
  assign n33598 = ~n11168 & n33597;
  assign n33599 = n11135 & n33598;
  assign n33600 = ~n11188 & n33599;
  assign n33601 = ~n14011 & n33600;
  assign n33602 = ~n14010 & n33601;
  assign n33603 = ~n12861 & n33602;
  assign n33604 = ~n12380 & n33603;
  assign n33605 = ~n12972 & n33604;
  assign n33606 = n14020 & n33605;
  assign n33607 = n13095 & n33606;
  assign n33608 = n14044 & n33607;
  assign n33609 = ~n33596 & ~n33608;
  assign n33610 = ~n33581 & n33609;
  assign n33611 = pi190 & ~n9717;
  assign n33612 = ~n9913 & n33611;
  assign n33613 = n9856 & n33612;
  assign n33614 = ~n9929 & n33613;
  assign n33615 = ~n13824 & n33614;
  assign n33616 = ~n13823 & n33615;
  assign n33617 = ~n11266 & n33616;
  assign n33618 = ~n12861 & n33617;
  assign n33619 = ~n11588 & n33618;
  assign n33620 = ~n12973 & n33619;
  assign n33621 = n13054 & n33620;
  assign n33622 = n13095 & n33621;
  assign n33623 = n13858 & n33622;
  assign n33624 = pi174 & ~n8574;
  assign n33625 = n11377 & n33624;
  assign n33626 = n9942 & n33625;
  assign n33627 = ~n8834 & n33626;
  assign n33628 = ~n10002 & n33627;
  assign n33629 = ~n13097 & n33628;
  assign n33630 = ~n13096 & n33629;
  assign n33631 = ~n11297 & n33630;
  assign n33632 = ~n12861 & n33631;
  assign n33633 = ~n12240 & n33632;
  assign n33634 = ~n12973 & n33633;
  assign n33635 = n13109 & n33634;
  assign n33636 = n13095 & n33635;
  assign n33637 = n13134 & n33636;
  assign n33638 = ~n33623 & ~n33637;
  assign n33639 = pi126 & ~n5627;
  assign n33640 = n5687 & n33639;
  assign n33641 = n13580 & n33640;
  assign n33642 = ~n5808 & n33641;
  assign n33643 = ~n6056 & n33642;
  assign n33644 = ~n7073 & n33643;
  assign n33645 = ~n8179 & n33644;
  assign n33646 = ~n9344 & n33645;
  assign n33647 = ~n13517 & n33646;
  assign n33648 = ~n13516 & n33647;
  assign n33649 = ~n10594 & n33648;
  assign n33650 = ~n12861 & n33649;
  assign n33651 = ~n12005 & n33650;
  assign n33652 = ~n13515 & n33651;
  assign n33653 = n13532 & n33652;
  assign n33654 = n13514 & n33653;
  assign n33655 = n13557 & n33654;
  assign n33656 = pi222 & ~n12671;
  assign n33657 = ~n12811 & n33656;
  assign n33658 = n13912 & n33657;
  assign n33659 = ~n12902 & n33658;
  assign n33660 = ~n13908 & n33659;
  assign n33661 = ~n12861 & n33660;
  assign n33662 = ~n12860 & n33661;
  assign n33663 = n12952 & n33662;
  assign n33664 = n13919 & n33663;
  assign n33665 = n14008 & n33664;
  assign n33666 = ~n33655 & ~n33665;
  assign n33667 = n33638 & n33666;
  assign n33668 = n13408 & n28569;
  assign n33669 = ~n3940 & n33668;
  assign n33670 = ~n4001 & n33669;
  assign n33671 = ~n5043 & n33670;
  assign n33672 = ~n5943 & n33671;
  assign n33673 = ~n6951 & n33672;
  assign n33674 = ~n8037 & n33673;
  assign n33675 = ~n9200 & n33674;
  assign n33676 = ~n13348 & n33675;
  assign n33677 = ~n13347 & n33676;
  assign n33678 = ~n10445 & n33677;
  assign n33679 = ~n12861 & n33678;
  assign n33680 = ~n11846 & n33679;
  assign n33681 = ~n13346 & n33680;
  assign n33682 = n13367 & n33681;
  assign n33683 = n13345 & n33682;
  assign n33684 = n13392 & n33683;
  assign n33685 = n13319 & n26369;
  assign n33686 = ~n3066 & n33685;
  assign n33687 = ~n3983 & n33686;
  assign n33688 = ~n4003 & n33687;
  assign n33689 = ~n4024 & n33688;
  assign n33690 = ~n4999 & n33689;
  assign n33691 = ~n5827 & n33690;
  assign n33692 = ~n6893 & n33691;
  assign n33693 = ~n7890 & n33692;
  assign n33694 = ~n9131 & n33693;
  assign n33695 = ~n13144 & n33694;
  assign n33696 = ~n13143 & n33695;
  assign n33697 = ~n10278 & n33696;
  assign n33698 = ~n13142 & n33697;
  assign n33699 = ~n11662 & n33698;
  assign n33700 = ~n13141 & n33699;
  assign n33701 = n13165 & n33700;
  assign n33702 = n13140 & n33701;
  assign n33703 = n13190 & n33702;
  assign n33704 = ~n33684 & ~n33703;
  assign n33705 = ~n12861 & n30988;
  assign n33706 = ~n12471 & n33705;
  assign n33707 = ~n12972 & n33706;
  assign n33708 = n14020 & n33707;
  assign n33709 = n13095 & n33708;
  assign n33710 = n14072 & n33709;
  assign n33711 = n13494 & n28602;
  assign n33712 = ~n4817 & n33711;
  assign n33713 = ~n4902 & n33712;
  assign n33714 = ~n6001 & n33713;
  assign n33715 = ~n7014 & n33714;
  assign n33716 = ~n8114 & n33715;
  assign n33717 = ~n9276 & n33716;
  assign n33718 = ~n13438 & n33717;
  assign n33719 = ~n13437 & n33718;
  assign n33720 = ~n10523 & n33719;
  assign n33721 = ~n12861 & n33720;
  assign n33722 = ~n11928 & n33721;
  assign n33723 = ~n13436 & n33722;
  assign n33724 = n13453 & n33723;
  assign n33725 = n13435 & n33724;
  assign n33726 = n13478 & n33725;
  assign n33727 = ~n33710 & ~n33726;
  assign n33728 = n33704 & n33727;
  assign n33729 = n33667 & n33728;
  assign n33730 = n33610 & n33729;
  assign po127 = ~n33574 | ~n33730;
  assign n33732 = n8485 & n31385;
  assign n33733 = ~n8834 & n33732;
  assign n33734 = ~n10002 & n33733;
  assign n33735 = ~n14747 & n33734;
  assign n33736 = ~n14746 & n33735;
  assign n33737 = ~n11297 & n33736;
  assign n33738 = ~n12240 & n33737;
  assign n33739 = ~n14467 & n33738;
  assign n33740 = ~n14466 & n33739;
  assign n33741 = n14574 & n33740;
  assign n33742 = n14760 & n33741;
  assign n33743 = n14764 & n33742;
  assign n33744 = n14745 & n33743;
  assign n33745 = n14787 & n33744;
  assign n33746 = ~n9913 & n26636;
  assign n33747 = n9794 & n33746;
  assign n33748 = ~n9929 & n33747;
  assign n33749 = ~n15497 & n33748;
  assign n33750 = ~n15496 & n33749;
  assign n33751 = ~n11266 & n33750;
  assign n33752 = ~n11588 & n33751;
  assign n33753 = ~n14467 & n33752;
  assign n33754 = ~n14466 & n33753;
  assign n33755 = n14574 & n33754;
  assign n33756 = n15508 & n33755;
  assign n33757 = n15512 & n33756;
  assign n33758 = n15495 & n33757;
  assign n33759 = n15535 & n33758;
  assign n33760 = ~n33745 & ~n33759;
  assign n33761 = pi231 & ~n14416;
  assign n33762 = n15890 & n33761;
  assign n33763 = ~n14519 & n33762;
  assign n33764 = ~n15742 & n33763;
  assign n33765 = ~n14467 & n33764;
  assign n33766 = ~n14466 & n33765;
  assign n33767 = n14574 & n33766;
  assign n33768 = ~n14577 & n33767;
  assign n33769 = n15756 & n33768;
  assign n33770 = n14457 & n33769;
  assign n33771 = n15854 & n33770;
  assign n33772 = ~n1205 & n31112;
  assign n33773 = ~n1203 & n33772;
  assign n33774 = ~n1238 & n33773;
  assign n33775 = n781 & n33774;
  assign n33776 = ~n1372 & n33775;
  assign n33777 = ~n2243 & n33776;
  assign n33778 = ~n3104 & n33777;
  assign n33779 = ~n3971 & n33778;
  assign n33780 = ~n4003 & n33779;
  assign n33781 = ~n4872 & n33780;
  assign n33782 = ~n5801 & n33781;
  assign n33783 = ~n6739 & n33782;
  assign n33784 = ~n7807 & n33783;
  assign n33785 = ~n8989 & n33784;
  assign n33786 = ~n10273 & n33785;
  assign n33787 = ~n14857 & n33786;
  assign n33788 = ~n14856 & n33787;
  assign n33789 = ~n11499 & n33788;
  assign n33790 = ~n13076 & n33789;
  assign n33791 = ~n14855 & n33790;
  assign n33792 = ~n14854 & n33791;
  assign n33793 = n14879 & n33792;
  assign n33794 = n14882 & n33793;
  assign n33795 = n14886 & n33794;
  assign n33796 = n14853 & n33795;
  assign n33797 = n14909 & n33796;
  assign n33798 = ~n33771 & ~n33797;
  assign n33799 = n33760 & n33798;
  assign n33800 = ~n12471 & n28799;
  assign n33801 = ~n14467 & n33800;
  assign n33802 = ~n14466 & n33801;
  assign n33803 = n14574 & n33802;
  assign n33804 = n15599 & n33803;
  assign n33805 = n15595 & n33804;
  assign n33806 = n15593 & n33805;
  assign n33807 = n15615 & n33806;
  assign n33808 = ~n12121 & n31081;
  assign n33809 = ~n14467 & n33808;
  assign n33810 = ~n13726 & n33809;
  assign n33811 = n14737 & n33810;
  assign n33812 = n15417 & n33811;
  assign n33813 = n15407 & n33812;
  assign n33814 = ~n11611 & n31096;
  assign n33815 = ~n14467 & n33814;
  assign n33816 = ~n13820 & n33815;
  assign n33817 = ~n14454 & n33816;
  assign n33818 = ~n14455 & n33817;
  assign n33819 = n14738 & n33818;
  assign n33820 = n14730 & n33819;
  assign n33821 = n14723 & n33820;
  assign n33822 = ~n33813 & ~n33821;
  assign n33823 = ~n33807 & n33822;
  assign n33824 = ~n13407 & n31142;
  assign n33825 = ~n14467 & n33824;
  assign n33826 = ~n15067 & n33825;
  assign n33827 = n15074 & n33826;
  assign n33828 = ~n13318 & n31146;
  assign n33829 = ~n14974 & n33828;
  assign n33830 = n14979 & n33829;
  assign n33831 = pi255 & ~n501;
  assign n33832 = n12872 & n33831;
  assign n33833 = n15973 & n33832;
  assign n33834 = n15980 & n33833;
  assign n33835 = n15972 & n33834;
  assign n33836 = n16005 & n33835;
  assign n33837 = ~n1172 & n33836;
  assign n33838 = ~n996 & n33837;
  assign n33839 = ~n2306 & n33838;
  assign n33840 = ~n500 & n33839;
  assign n33841 = n16011 & n33840;
  assign n33842 = n16014 & n33841;
  assign n33843 = n16017 & n33842;
  assign n33844 = n16038 & n33843;
  assign n33845 = n15963 & n33844;
  assign n33846 = n15954 & n33845;
  assign n33847 = ~n7236 & n33846;
  assign n33848 = ~n6137 & n33847;
  assign n33849 = n6193 & n33848;
  assign n33850 = n6134 & n33849;
  assign n33851 = ~n8867 & n33850;
  assign n33852 = ~n7235 & n33851;
  assign n33853 = n7296 & n33852;
  assign n33854 = n7231 & n33853;
  assign n33855 = ~n10027 & n33854;
  assign n33856 = ~n8866 & n33855;
  assign n33857 = n8898 & n33856;
  assign n33858 = n8863 & n33857;
  assign n33859 = pi247 & ~n501;
  assign n33860 = n12872 & n33859;
  assign n33861 = n15973 & n33860;
  assign n33862 = n16069 & n33861;
  assign n33863 = n16063 & n33862;
  assign n33864 = n16088 & n33863;
  assign n33865 = ~n1172 & n33864;
  assign n33866 = ~n996 & n33865;
  assign n33867 = ~n2306 & n33866;
  assign n33868 = ~n500 & n33867;
  assign n33869 = n16094 & n33868;
  assign n33870 = n16016 & n33869;
  assign n33871 = n16054 & n33870;
  assign n33872 = n16113 & n33871;
  assign n33873 = n16184 & n33872;
  assign n33874 = n16048 & n33873;
  assign n33875 = ~n7236 & n33874;
  assign n33876 = ~n6137 & n33875;
  assign n33877 = n6193 & n33876;
  assign n33878 = n6134 & n33877;
  assign n33879 = ~n8867 & n33878;
  assign n33880 = ~n7235 & n33879;
  assign n33881 = n7296 & n33880;
  assign n33882 = n7231 & n33881;
  assign n33883 = ~n10027 & n33882;
  assign n33884 = ~n8866 & n33883;
  assign n33885 = n8898 & n33884;
  assign n33886 = n8863 & n33885;
  assign n33887 = ~n33858 & ~n33886;
  assign n33888 = ~n10788 & ~n33887;
  assign n33889 = ~n10026 & n33888;
  assign n33890 = n10072 & n33889;
  assign n33891 = n10021 & n33890;
  assign n33892 = ~n33830 & ~n33891;
  assign n33893 = ~n33827 & n33892;
  assign n33894 = ~n13579 & n31231;
  assign n33895 = ~n14467 & n33894;
  assign n33896 = n14574 & n33895;
  assign n33897 = ~n15270 & n33896;
  assign n33898 = n15276 & n33897;
  assign n33899 = n15269 & n33898;
  assign n33900 = ~n13493 & n31226;
  assign n33901 = ~n14467 & n33900;
  assign n33902 = ~n14573 & n33901;
  assign n33903 = ~n15156 & n33902;
  assign n33904 = n15166 & n33903;
  assign n33905 = ~n33899 & ~n33904;
  assign n33906 = n33893 & n33905;
  assign n33907 = ~n12181 & n31088;
  assign n33908 = ~n14467 & n33907;
  assign n33909 = ~n13764 & n33908;
  assign n33910 = ~n14455 & n33909;
  assign n33911 = n14737 & n33910;
  assign n33912 = n15463 & n33911;
  assign n33913 = n15452 & n33912;
  assign n33914 = ~n11551 & n31103;
  assign n33915 = ~n14467 & n33914;
  assign n33916 = ~n13906 & n33915;
  assign n33917 = ~n14452 & n33916;
  assign n33918 = n14456 & n33917;
  assign n33919 = n15571 & n33918;
  assign n33920 = n15585 & n33919;
  assign n33921 = ~n33913 & ~n33920;
  assign n33922 = n33906 & n33921;
  assign n33923 = n33823 & n33922;
  assign n33924 = n33799 & n33923;
  assign n33925 = ~n4401 & n31254;
  assign n33926 = n4490 & n33925;
  assign n33927 = ~n4817 & n33926;
  assign n33928 = ~n4902 & n33927;
  assign n33929 = ~n6001 & n33928;
  assign n33930 = ~n7014 & n33929;
  assign n33931 = ~n8114 & n33930;
  assign n33932 = ~n9276 & n33931;
  assign n33933 = ~n15107 & n33932;
  assign n33934 = ~n15106 & n33933;
  assign n33935 = ~n10523 & n33934;
  assign n33936 = ~n11928 & n33935;
  assign n33937 = ~n14467 & n33936;
  assign n33938 = ~n14573 & n33937;
  assign n33939 = n15122 & n33938;
  assign n33940 = n15125 & n33939;
  assign n33941 = n15129 & n33940;
  assign n33942 = n15105 & n33941;
  assign n33943 = n15152 & n33942;
  assign n33944 = pi239 & ~n14568;
  assign n33945 = ~n14520 & n33944;
  assign n33946 = ~n14467 & n33945;
  assign n33947 = ~n14466 & n33946;
  assign n33948 = n14574 & n33947;
  assign n33949 = ~n14465 & n33948;
  assign n33950 = n14581 & n33949;
  assign n33951 = n14457 & n33950;
  assign n33952 = n14715 & n33951;
  assign n33953 = n1738 & n31334;
  assign n33954 = ~n1735 & n33953;
  assign n33955 = ~n1521 & n33954;
  assign n33956 = ~n1556 & n33955;
  assign n33957 = ~n1587 & n33956;
  assign n33958 = ~n2242 & n33957;
  assign n33959 = ~n3095 & n33958;
  assign n33960 = ~n3997 & n33959;
  assign n33961 = ~n4003 & n33960;
  assign n33962 = ~n4837 & n33961;
  assign n33963 = ~n5822 & n33962;
  assign n33964 = ~n6820 & n33963;
  assign n33965 = ~n7785 & n33964;
  assign n33966 = ~n9027 & n33965;
  assign n33967 = ~n10245 & n33966;
  assign n33968 = ~n14919 & n33967;
  assign n33969 = ~n14918 & n33968;
  assign n33970 = ~n11536 & n33969;
  assign n33971 = ~n13036 & n33970;
  assign n33972 = ~n14917 & n33971;
  assign n33973 = ~n14916 & n33972;
  assign n33974 = n14940 & n33973;
  assign n33975 = n14943 & n33974;
  assign n33976 = n14947 & n33975;
  assign n33977 = n14915 & n33976;
  assign n33978 = n14970 & n33977;
  assign n33979 = ~n33952 & ~n33978;
  assign n33980 = ~n33943 & n33979;
  assign n33981 = ~n14467 & n31309;
  assign n33982 = ~n14466 & n33981;
  assign n33983 = n14574 & n33982;
  assign n33984 = n15859 & n33983;
  assign n33985 = n15862 & n33984;
  assign n33986 = n15595 & n33985;
  assign n33987 = n15885 & n33986;
  assign n33988 = n4103 & n31361;
  assign n33989 = ~n3940 & n33988;
  assign n33990 = ~n4001 & n33989;
  assign n33991 = ~n5043 & n33990;
  assign n33992 = ~n5943 & n33991;
  assign n33993 = ~n6951 & n33992;
  assign n33994 = ~n8037 & n33993;
  assign n33995 = ~n9200 & n33994;
  assign n33996 = ~n15012 & n33995;
  assign n33997 = ~n15011 & n33996;
  assign n33998 = ~n10445 & n33997;
  assign n33999 = ~n11846 & n33998;
  assign n34000 = ~n14467 & n33999;
  assign n34001 = ~n15010 & n34000;
  assign n34002 = n15030 & n34001;
  assign n34003 = n15033 & n34002;
  assign n34004 = n15037 & n34003;
  assign n34005 = n15009 & n34004;
  assign n34006 = n15060 & n34005;
  assign n34007 = ~n33987 & ~n34006;
  assign n34008 = n15386 & n31316;
  assign n34009 = ~n6784 & n34008;
  assign n34010 = ~n7158 & n34009;
  assign n34011 = ~n8250 & n34010;
  assign n34012 = ~n9414 & n34011;
  assign n34013 = ~n15287 & n34012;
  assign n34014 = ~n15286 & n34013;
  assign n34015 = ~n10667 & n34014;
  assign n34016 = ~n12083 & n34015;
  assign n34017 = ~n14467 & n34016;
  assign n34018 = ~n14466 & n34017;
  assign n34019 = n14574 & n34018;
  assign n34020 = n15302 & n34019;
  assign n34021 = n15306 & n34020;
  assign n34022 = n15285 & n34021;
  assign n34023 = n15329 & n34022;
  assign n34024 = pi151 & ~n7663;
  assign n34025 = n15424 & n34024;
  assign n34026 = ~n7869 & n34025;
  assign n34027 = ~n8346 & n34026;
  assign n34028 = ~n9485 & n34027;
  assign n34029 = ~n15345 & n34028;
  assign n34030 = ~n15344 & n34029;
  assign n34031 = ~n10741 & n34030;
  assign n34032 = ~n12158 & n34031;
  assign n34033 = ~n14467 & n34032;
  assign n34034 = ~n14466 & n34033;
  assign n34035 = n14574 & n34034;
  assign n34036 = n15357 & n34035;
  assign n34037 = n15361 & n34036;
  assign n34038 = n15343 & n34037;
  assign n34039 = n15384 & n34038;
  assign n34040 = ~n34023 & ~n34039;
  assign n34041 = n34007 & n34040;
  assign n34042 = n3846 & n31415;
  assign n34043 = ~n3066 & n34042;
  assign n34044 = ~n3983 & n34043;
  assign n34045 = ~n4003 & n34044;
  assign n34046 = ~n4024 & n34045;
  assign n34047 = ~n4999 & n34046;
  assign n34048 = ~n5827 & n34047;
  assign n34049 = ~n6893 & n34048;
  assign n34050 = ~n7890 & n34049;
  assign n34051 = ~n9131 & n34050;
  assign n34052 = ~n14797 & n34051;
  assign n34053 = ~n14796 & n34052;
  assign n34054 = ~n10278 & n34053;
  assign n34055 = ~n11662 & n34054;
  assign n34056 = ~n14795 & n34055;
  assign n34057 = ~n14794 & n34056;
  assign n34058 = n14817 & n34057;
  assign n34059 = n14820 & n34058;
  assign n34060 = n14824 & n34059;
  assign n34061 = n14793 & n34060;
  assign n34062 = n14847 & n34061;
  assign n34063 = pi199 & ~n11168;
  assign n34064 = n15698 & n34063;
  assign n34065 = ~n11188 & n34064;
  assign n34066 = ~n15620 & n34065;
  assign n34067 = ~n15619 & n34066;
  assign n34068 = ~n12380 & n34067;
  assign n34069 = ~n14467 & n34068;
  assign n34070 = ~n14466 & n34069;
  assign n34071 = n14574 & n34070;
  assign n34072 = n15629 & n34071;
  assign n34073 = n15633 & n34072;
  assign n34074 = n15595 & n34073;
  assign n34075 = n15656 & n34074;
  assign n34076 = ~n34062 & ~n34075;
  assign n34077 = pi215 & ~n12841;
  assign n34078 = n12775 & n34077;
  assign n34079 = ~n12902 & n34078;
  assign n34080 = ~n15659 & n34079;
  assign n34081 = ~n15658 & n34080;
  assign n34082 = ~n14467 & n34081;
  assign n34083 = ~n14466 & n34082;
  assign n34084 = n14574 & n34083;
  assign n34085 = n15666 & n34084;
  assign n34086 = n15669 & n34085;
  assign n34087 = n15595 & n34086;
  assign n34088 = n15692 & n34087;
  assign n34089 = n15247 & n31435;
  assign n34090 = ~n5808 & n34089;
  assign n34091 = ~n6056 & n34090;
  assign n34092 = ~n7073 & n34091;
  assign n34093 = ~n8179 & n34092;
  assign n34094 = ~n9344 & n34093;
  assign n34095 = ~n15195 & n34094;
  assign n34096 = ~n15194 & n34095;
  assign n34097 = ~n10594 & n34096;
  assign n34098 = ~n12005 & n34097;
  assign n34099 = ~n14467 & n34098;
  assign n34100 = ~n14572 & n34099;
  assign n34101 = n15208 & n34100;
  assign n34102 = n15211 & n34101;
  assign n34103 = n15215 & n34102;
  assign n34104 = n15193 & n34103;
  assign n34105 = n15238 & n34104;
  assign n34106 = ~n34088 & ~n34105;
  assign n34107 = n34076 & n34106;
  assign n34108 = n34041 & n34107;
  assign n34109 = n33980 & n34108;
  assign po128 = ~n33924 | ~n34109;
  assign n34111 = pi104 & ~n4401;
  assign n34112 = n13494 & n34111;
  assign n34113 = ~n4817 & n34112;
  assign n34114 = ~n4902 & n34113;
  assign n34115 = ~n6001 & n34114;
  assign n34116 = ~n7014 & n34115;
  assign n34117 = ~n8114 & n34116;
  assign n34118 = ~n9276 & n34117;
  assign n34119 = ~n15107 & n34118;
  assign n34120 = ~n15106 & n34119;
  assign n34121 = ~n10523 & n34120;
  assign n34122 = ~n11928 & n34121;
  assign n34123 = ~n14467 & n34122;
  assign n34124 = ~n14573 & n34123;
  assign n34125 = n15122 & n34124;
  assign n34126 = n15125 & n34125;
  assign n34127 = n15129 & n34126;
  assign n34128 = n15105 & n34127;
  assign n34129 = n15152 & n34128;
  assign n34130 = n15386 & n27007;
  assign n34131 = ~n6784 & n34130;
  assign n34132 = ~n7158 & n34131;
  assign n34133 = ~n8250 & n34132;
  assign n34134 = ~n9414 & n34133;
  assign n34135 = ~n15287 & n34134;
  assign n34136 = ~n15286 & n34135;
  assign n34137 = ~n10667 & n34136;
  assign n34138 = ~n12083 & n34137;
  assign n34139 = ~n14467 & n34138;
  assign n34140 = ~n14466 & n34139;
  assign n34141 = n14574 & n34140;
  assign n34142 = n15302 & n34141;
  assign n34143 = n15306 & n34142;
  assign n34144 = n15285 & n34143;
  assign n34145 = n15329 & n34144;
  assign n34146 = ~n34129 & ~n34145;
  assign n34147 = n13408 & n26787;
  assign n34148 = ~n3940 & n34147;
  assign n34149 = ~n4001 & n34148;
  assign n34150 = ~n5043 & n34149;
  assign n34151 = ~n5943 & n34150;
  assign n34152 = ~n6951 & n34151;
  assign n34153 = ~n8037 & n34152;
  assign n34154 = ~n9200 & n34153;
  assign n34155 = ~n15012 & n34154;
  assign n34156 = ~n15011 & n34155;
  assign n34157 = ~n10445 & n34156;
  assign n34158 = ~n11846 & n34157;
  assign n34159 = ~n14467 & n34158;
  assign n34160 = ~n15010 & n34159;
  assign n34161 = n15030 & n34160;
  assign n34162 = n15033 & n34161;
  assign n34163 = n15037 & n34162;
  assign n34164 = n15009 & n34163;
  assign n34165 = n15060 & n34164;
  assign n34166 = pi184 & ~n9913;
  assign n34167 = n15548 & n34166;
  assign n34168 = ~n9929 & n34167;
  assign n34169 = ~n15497 & n34168;
  assign n34170 = ~n15496 & n34169;
  assign n34171 = ~n11266 & n34170;
  assign n34172 = ~n11588 & n34171;
  assign n34173 = ~n14467 & n34172;
  assign n34174 = ~n14466 & n34173;
  assign n34175 = n14574 & n34174;
  assign n34176 = n15508 & n34175;
  assign n34177 = n15512 & n34176;
  assign n34178 = n15495 & n34177;
  assign n34179 = n15535 & n34178;
  assign n34180 = ~n34165 & ~n34179;
  assign n34181 = n34146 & n34180;
  assign n34182 = ~n12471 & n29169;
  assign n34183 = ~n14467 & n34182;
  assign n34184 = ~n14466 & n34183;
  assign n34185 = n14574 & n34184;
  assign n34186 = n15599 & n34185;
  assign n34187 = n15595 & n34186;
  assign n34188 = n15593 & n34187;
  assign n34189 = n15615 & n34188;
  assign n34190 = ~n11611 & n31479;
  assign n34191 = ~n14467 & n34190;
  assign n34192 = ~n13820 & n34191;
  assign n34193 = ~n14454 & n34192;
  assign n34194 = ~n14455 & n34193;
  assign n34195 = n14738 & n34194;
  assign n34196 = n14730 & n34195;
  assign n34197 = n14723 & n34196;
  assign n34198 = ~n11551 & n31457;
  assign n34199 = ~n14467 & n34198;
  assign n34200 = ~n13906 & n34199;
  assign n34201 = ~n14452 & n34200;
  assign n34202 = n14456 & n34201;
  assign n34203 = n15571 & n34202;
  assign n34204 = n15585 & n34203;
  assign n34205 = ~n34197 & ~n34204;
  assign n34206 = ~n34189 & n34205;
  assign n34207 = ~n13579 & n31501;
  assign n34208 = ~n14467 & n34207;
  assign n34209 = n14574 & n34208;
  assign n34210 = ~n15270 & n34209;
  assign n34211 = n15276 & n34210;
  assign n34212 = n15269 & n34211;
  assign n34213 = pi256 & ~n501;
  assign n34214 = n12872 & n34213;
  assign n34215 = n15973 & n34214;
  assign n34216 = n15980 & n34215;
  assign n34217 = n15972 & n34216;
  assign n34218 = n16005 & n34217;
  assign n34219 = ~n1172 & n34218;
  assign n34220 = ~n996 & n34219;
  assign n34221 = ~n2306 & n34220;
  assign n34222 = ~n500 & n34221;
  assign n34223 = n16011 & n34222;
  assign n34224 = n16014 & n34223;
  assign n34225 = n16017 & n34224;
  assign n34226 = n16038 & n34225;
  assign n34227 = n15963 & n34226;
  assign n34228 = n15954 & n34227;
  assign n34229 = ~n7236 & n34228;
  assign n34230 = ~n6137 & n34229;
  assign n34231 = n6193 & n34230;
  assign n34232 = n6134 & n34231;
  assign n34233 = ~n8867 & n34232;
  assign n34234 = ~n7235 & n34233;
  assign n34235 = n7296 & n34234;
  assign n34236 = n7231 & n34235;
  assign n34237 = ~n10027 & n34236;
  assign n34238 = ~n8866 & n34237;
  assign n34239 = n8898 & n34238;
  assign n34240 = n8863 & n34239;
  assign n34241 = pi248 & ~n501;
  assign n34242 = n12872 & n34241;
  assign n34243 = n15973 & n34242;
  assign n34244 = n16069 & n34243;
  assign n34245 = n16063 & n34244;
  assign n34246 = n16088 & n34245;
  assign n34247 = ~n1172 & n34246;
  assign n34248 = ~n996 & n34247;
  assign n34249 = ~n2306 & n34248;
  assign n34250 = ~n500 & n34249;
  assign n34251 = n16094 & n34250;
  assign n34252 = n16016 & n34251;
  assign n34253 = n16054 & n34252;
  assign n34254 = n16113 & n34253;
  assign n34255 = n16184 & n34254;
  assign n34256 = n16048 & n34255;
  assign n34257 = ~n7236 & n34256;
  assign n34258 = ~n6137 & n34257;
  assign n34259 = n6193 & n34258;
  assign n34260 = n6134 & n34259;
  assign n34261 = ~n8867 & n34260;
  assign n34262 = ~n7235 & n34261;
  assign n34263 = n7296 & n34262;
  assign n34264 = n7231 & n34263;
  assign n34265 = ~n10027 & n34264;
  assign n34266 = ~n8866 & n34265;
  assign n34267 = n8898 & n34266;
  assign n34268 = n8863 & n34267;
  assign n34269 = ~n34240 & ~n34268;
  assign n34270 = ~n10788 & ~n34269;
  assign n34271 = ~n10026 & n34270;
  assign n34272 = n10072 & n34271;
  assign n34273 = n10021 & n34272;
  assign n34274 = ~n13318 & n31506;
  assign n34275 = ~n14974 & n34274;
  assign n34276 = n14979 & n34275;
  assign n34277 = ~n34273 & ~n34276;
  assign n34278 = ~n34212 & n34277;
  assign n34279 = ~n13407 & n31567;
  assign n34280 = ~n14467 & n34279;
  assign n34281 = ~n15067 & n34280;
  assign n34282 = n15074 & n34281;
  assign n34283 = ~n13493 & n31571;
  assign n34284 = ~n14467 & n34283;
  assign n34285 = ~n14573 & n34284;
  assign n34286 = ~n15156 & n34285;
  assign n34287 = n15166 & n34286;
  assign n34288 = ~n34282 & ~n34287;
  assign n34289 = n34278 & n34288;
  assign n34290 = ~n12121 & n31464;
  assign n34291 = ~n14467 & n34290;
  assign n34292 = ~n13726 & n34291;
  assign n34293 = n14737 & n34292;
  assign n34294 = n15417 & n34293;
  assign n34295 = n15407 & n34294;
  assign n34296 = ~n12181 & n31472;
  assign n34297 = ~n14467 & n34296;
  assign n34298 = ~n13764 & n34297;
  assign n34299 = ~n14455 & n34298;
  assign n34300 = n14737 & n34299;
  assign n34301 = n15463 & n34300;
  assign n34302 = n15452 & n34301;
  assign n34303 = ~n34295 & ~n34302;
  assign n34304 = n34289 & n34303;
  assign n34305 = n34206 & n34304;
  assign n34306 = n34181 & n34305;
  assign n34307 = ~n14467 & n31675;
  assign n34308 = ~n14466 & n34307;
  assign n34309 = n14574 & n34308;
  assign n34310 = n15859 & n34309;
  assign n34311 = n15862 & n34310;
  assign n34312 = n15595 & n34311;
  assign n34313 = n15885 & n34312;
  assign n34314 = pi240 & ~n14568;
  assign n34315 = ~n14520 & n34314;
  assign n34316 = ~n14467 & n34315;
  assign n34317 = ~n14466 & n34316;
  assign n34318 = n14574 & n34317;
  assign n34319 = ~n14465 & n34318;
  assign n34320 = n14581 & n34319;
  assign n34321 = n14457 & n34320;
  assign n34322 = n14715 & n34321;
  assign n34323 = pi056 & ~n1740;
  assign n34324 = n13259 & n34323;
  assign n34325 = ~n2242 & n34324;
  assign n34326 = ~n3095 & n34325;
  assign n34327 = ~n3997 & n34326;
  assign n34328 = ~n4003 & n34327;
  assign n34329 = ~n4837 & n34328;
  assign n34330 = ~n5822 & n34329;
  assign n34331 = ~n6820 & n34330;
  assign n34332 = ~n7785 & n34331;
  assign n34333 = ~n9027 & n34332;
  assign n34334 = ~n10245 & n34333;
  assign n34335 = ~n14919 & n34334;
  assign n34336 = ~n14918 & n34335;
  assign n34337 = ~n11536 & n34336;
  assign n34338 = ~n13036 & n34337;
  assign n34339 = ~n14917 & n34338;
  assign n34340 = ~n14916 & n34339;
  assign n34341 = n14940 & n34340;
  assign n34342 = n14943 & n34341;
  assign n34343 = n14947 & n34342;
  assign n34344 = n14915 & n34343;
  assign n34345 = n14970 & n34344;
  assign n34346 = ~n34322 & ~n34345;
  assign n34347 = ~n34313 & n34346;
  assign n34348 = n14749 & n31592;
  assign n34349 = ~n8834 & n34348;
  assign n34350 = ~n10002 & n34349;
  assign n34351 = ~n14747 & n34350;
  assign n34352 = ~n14746 & n34351;
  assign n34353 = ~n11297 & n34352;
  assign n34354 = ~n12240 & n34353;
  assign n34355 = ~n14467 & n34354;
  assign n34356 = ~n14466 & n34355;
  assign n34357 = n14574 & n34356;
  assign n34358 = n14760 & n34357;
  assign n34359 = n14764 & n34358;
  assign n34360 = n14745 & n34359;
  assign n34361 = n14787 & n34360;
  assign n34362 = n15424 & n23403;
  assign n34363 = ~n7869 & n34362;
  assign n34364 = ~n8346 & n34363;
  assign n34365 = ~n9485 & n34364;
  assign n34366 = ~n15345 & n34365;
  assign n34367 = ~n15344 & n34366;
  assign n34368 = ~n10741 & n34367;
  assign n34369 = ~n12158 & n34368;
  assign n34370 = ~n14467 & n34369;
  assign n34371 = ~n14466 & n34370;
  assign n34372 = n14574 & n34371;
  assign n34373 = n15357 & n34372;
  assign n34374 = n15361 & n34373;
  assign n34375 = n15343 & n34374;
  assign n34376 = n15384 & n34375;
  assign n34377 = ~n34361 & ~n34376;
  assign n34378 = n15247 & n31760;
  assign n34379 = ~n5808 & n34378;
  assign n34380 = ~n6056 & n34379;
  assign n34381 = ~n7073 & n34380;
  assign n34382 = ~n8179 & n34381;
  assign n34383 = ~n9344 & n34382;
  assign n34384 = ~n15195 & n34383;
  assign n34385 = ~n15194 & n34384;
  assign n34386 = ~n10594 & n34385;
  assign n34387 = ~n12005 & n34386;
  assign n34388 = ~n14467 & n34387;
  assign n34389 = ~n14572 & n34388;
  assign n34390 = n15208 & n34389;
  assign n34391 = n15211 & n34390;
  assign n34392 = n15215 & n34391;
  assign n34393 = n15193 & n34392;
  assign n34394 = n15238 & n34393;
  assign n34395 = pi200 & ~n11168;
  assign n34396 = n15698 & n34395;
  assign n34397 = ~n11188 & n34396;
  assign n34398 = ~n15620 & n34397;
  assign n34399 = ~n15619 & n34398;
  assign n34400 = ~n12380 & n34399;
  assign n34401 = ~n14467 & n34400;
  assign n34402 = ~n14466 & n34401;
  assign n34403 = n14574 & n34402;
  assign n34404 = n15629 & n34403;
  assign n34405 = n15633 & n34404;
  assign n34406 = n15595 & n34405;
  assign n34407 = n15656 & n34406;
  assign n34408 = ~n34394 & ~n34407;
  assign n34409 = n34377 & n34408;
  assign n34410 = pi216 & ~n12841;
  assign n34411 = n12775 & n34410;
  assign n34412 = ~n12902 & n34411;
  assign n34413 = ~n15659 & n34412;
  assign n34414 = ~n15658 & n34413;
  assign n34415 = ~n14467 & n34414;
  assign n34416 = ~n14466 & n34415;
  assign n34417 = n14574 & n34416;
  assign n34418 = n15666 & n34417;
  assign n34419 = n15669 & n34418;
  assign n34420 = n15595 & n34419;
  assign n34421 = n15692 & n34420;
  assign n34422 = pi232 & ~n14416;
  assign n34423 = n15890 & n34422;
  assign n34424 = ~n14519 & n34423;
  assign n34425 = ~n15742 & n34424;
  assign n34426 = ~n14467 & n34425;
  assign n34427 = ~n14466 & n34426;
  assign n34428 = n14574 & n34427;
  assign n34429 = ~n14577 & n34428;
  assign n34430 = n15756 & n34429;
  assign n34431 = n14457 & n34430;
  assign n34432 = n15854 & n34431;
  assign n34433 = ~n34421 & ~n34432;
  assign n34434 = n14858 & n26952;
  assign n34435 = ~n1372 & n34434;
  assign n34436 = ~n2243 & n34435;
  assign n34437 = ~n3104 & n34436;
  assign n34438 = ~n3971 & n34437;
  assign n34439 = ~n4003 & n34438;
  assign n34440 = ~n4872 & n34439;
  assign n34441 = ~n5801 & n34440;
  assign n34442 = ~n6739 & n34441;
  assign n34443 = ~n7807 & n34442;
  assign n34444 = ~n8989 & n34443;
  assign n34445 = ~n10273 & n34444;
  assign n34446 = ~n14857 & n34445;
  assign n34447 = ~n14856 & n34446;
  assign n34448 = ~n11499 & n34447;
  assign n34449 = ~n13076 & n34448;
  assign n34450 = ~n14855 & n34449;
  assign n34451 = ~n14854 & n34450;
  assign n34452 = n14879 & n34451;
  assign n34453 = n14882 & n34452;
  assign n34454 = n14886 & n34453;
  assign n34455 = n14853 & n34454;
  assign n34456 = n14909 & n34455;
  assign n34457 = n14981 & n21883;
  assign n34458 = ~n3066 & n34457;
  assign n34459 = ~n3983 & n34458;
  assign n34460 = ~n4003 & n34459;
  assign n34461 = ~n4024 & n34460;
  assign n34462 = ~n4999 & n34461;
  assign n34463 = ~n5827 & n34462;
  assign n34464 = ~n6893 & n34463;
  assign n34465 = ~n7890 & n34464;
  assign n34466 = ~n9131 & n34465;
  assign n34467 = ~n14797 & n34466;
  assign n34468 = ~n14796 & n34467;
  assign n34469 = ~n10278 & n34468;
  assign n34470 = ~n11662 & n34469;
  assign n34471 = ~n14795 & n34470;
  assign n34472 = ~n14794 & n34471;
  assign n34473 = n14817 & n34472;
  assign n34474 = n14820 & n34473;
  assign n34475 = n14824 & n34474;
  assign n34476 = n14793 & n34475;
  assign n34477 = n14847 & n34476;
  assign n34478 = ~n34456 & ~n34477;
  assign n34479 = n34433 & n34478;
  assign n34480 = n34409 & n34479;
  assign n34481 = n34347 & n34480;
  assign po129 = ~n34306 | ~n34481;
  assign n34483 = pi057 & ~n1740;
  assign n34484 = n13259 & n34483;
  assign n34485 = ~n2242 & n34484;
  assign n34486 = ~n3095 & n34485;
  assign n34487 = ~n3997 & n34486;
  assign n34488 = ~n4003 & n34487;
  assign n34489 = ~n4837 & n34488;
  assign n34490 = ~n5822 & n34489;
  assign n34491 = ~n6820 & n34490;
  assign n34492 = ~n7785 & n34491;
  assign n34493 = ~n9027 & n34492;
  assign n34494 = ~n10245 & n34493;
  assign n34495 = ~n14919 & n34494;
  assign n34496 = ~n14918 & n34495;
  assign n34497 = ~n11536 & n34496;
  assign n34498 = ~n13036 & n34497;
  assign n34499 = ~n14917 & n34498;
  assign n34500 = ~n14916 & n34499;
  assign n34501 = n14940 & n34500;
  assign n34502 = n14943 & n34501;
  assign n34503 = n14947 & n34502;
  assign n34504 = n14915 & n34503;
  assign n34505 = n14970 & n34504;
  assign n34506 = pi217 & ~n12841;
  assign n34507 = n12775 & n34506;
  assign n34508 = ~n12902 & n34507;
  assign n34509 = ~n15659 & n34508;
  assign n34510 = ~n15658 & n34509;
  assign n34511 = ~n14467 & n34510;
  assign n34512 = ~n14466 & n34511;
  assign n34513 = n14574 & n34512;
  assign n34514 = n15666 & n34513;
  assign n34515 = n15669 & n34514;
  assign n34516 = n15595 & n34515;
  assign n34517 = n15692 & n34516;
  assign n34518 = ~n34505 & ~n34517;
  assign n34519 = ~n14467 & n32017;
  assign n34520 = ~n14466 & n34519;
  assign n34521 = n14574 & n34520;
  assign n34522 = n15859 & n34521;
  assign n34523 = n15862 & n34522;
  assign n34524 = n15595 & n34523;
  assign n34525 = n15885 & n34524;
  assign n34526 = n14749 & n32003;
  assign n34527 = ~n8834 & n34526;
  assign n34528 = ~n10002 & n34527;
  assign n34529 = ~n14747 & n34528;
  assign n34530 = ~n14746 & n34529;
  assign n34531 = ~n11297 & n34530;
  assign n34532 = ~n12240 & n34531;
  assign n34533 = ~n14467 & n34532;
  assign n34534 = ~n14466 & n34533;
  assign n34535 = n14574 & n34534;
  assign n34536 = n14760 & n34535;
  assign n34537 = n14764 & n34536;
  assign n34538 = n14745 & n34537;
  assign n34539 = n14787 & n34538;
  assign n34540 = ~n34525 & ~n34539;
  assign n34541 = n34518 & n34540;
  assign n34542 = ~n11611 & n31782;
  assign n34543 = ~n14467 & n34542;
  assign n34544 = ~n13820 & n34543;
  assign n34545 = ~n14454 & n34544;
  assign n34546 = ~n14455 & n34545;
  assign n34547 = n14738 & n34546;
  assign n34548 = n14730 & n34547;
  assign n34549 = n14723 & n34548;
  assign n34550 = ~n12181 & n31797;
  assign n34551 = ~n14467 & n34550;
  assign n34552 = ~n13764 & n34551;
  assign n34553 = ~n14455 & n34552;
  assign n34554 = n14737 & n34553;
  assign n34555 = n15463 & n34554;
  assign n34556 = n15452 & n34555;
  assign n34557 = ~n11551 & n31804;
  assign n34558 = ~n14467 & n34557;
  assign n34559 = ~n13906 & n34558;
  assign n34560 = ~n14452 & n34559;
  assign n34561 = n14456 & n34560;
  assign n34562 = n15571 & n34561;
  assign n34563 = n15585 & n34562;
  assign n34564 = ~n34556 & ~n34563;
  assign n34565 = ~n34549 & n34564;
  assign n34566 = ~n13579 & n31905;
  assign n34567 = ~n14467 & n34566;
  assign n34568 = n14574 & n34567;
  assign n34569 = ~n15270 & n34568;
  assign n34570 = n15276 & n34569;
  assign n34571 = n15269 & n34570;
  assign n34572 = pi249 & ~n501;
  assign n34573 = n12872 & n34572;
  assign n34574 = n15973 & n34573;
  assign n34575 = n16069 & n34574;
  assign n34576 = n16063 & n34575;
  assign n34577 = n16088 & n34576;
  assign n34578 = ~n1172 & n34577;
  assign n34579 = ~n996 & n34578;
  assign n34580 = ~n2306 & n34579;
  assign n34581 = ~n500 & n34580;
  assign n34582 = n16094 & n34581;
  assign n34583 = n16016 & n34582;
  assign n34584 = n16054 & n34583;
  assign n34585 = n16113 & n34584;
  assign n34586 = n16184 & n34585;
  assign n34587 = n16048 & n34586;
  assign n34588 = ~n7236 & n34587;
  assign n34589 = ~n6137 & n34588;
  assign n34590 = n6193 & n34589;
  assign n34591 = n6134 & n34590;
  assign n34592 = ~n8867 & n34591;
  assign n34593 = ~n7235 & n34592;
  assign n34594 = n7296 & n34593;
  assign n34595 = n7231 & n34594;
  assign n34596 = ~n10027 & n34595;
  assign n34597 = ~n8866 & n34596;
  assign n34598 = n8898 & n34597;
  assign n34599 = n8863 & n34598;
  assign n34600 = pi257 & ~n501;
  assign n34601 = n12872 & n34600;
  assign n34602 = n15973 & n34601;
  assign n34603 = n15980 & n34602;
  assign n34604 = n15972 & n34603;
  assign n34605 = n16005 & n34604;
  assign n34606 = ~n1172 & n34605;
  assign n34607 = ~n996 & n34606;
  assign n34608 = ~n2306 & n34607;
  assign n34609 = ~n500 & n34608;
  assign n34610 = n16011 & n34609;
  assign n34611 = n16014 & n34610;
  assign n34612 = n16017 & n34611;
  assign n34613 = n16038 & n34612;
  assign n34614 = n15963 & n34613;
  assign n34615 = n15954 & n34614;
  assign n34616 = ~n7236 & n34615;
  assign n34617 = ~n6137 & n34616;
  assign n34618 = n6193 & n34617;
  assign n34619 = n6134 & n34618;
  assign n34620 = ~n8867 & n34619;
  assign n34621 = ~n7235 & n34620;
  assign n34622 = n7296 & n34621;
  assign n34623 = n7231 & n34622;
  assign n34624 = ~n10027 & n34623;
  assign n34625 = ~n8866 & n34624;
  assign n34626 = n8898 & n34625;
  assign n34627 = n8863 & n34626;
  assign n34628 = ~n34599 & ~n34627;
  assign n34629 = ~n10788 & ~n34628;
  assign n34630 = ~n10026 & n34629;
  assign n34631 = n10072 & n34630;
  assign n34632 = n10021 & n34631;
  assign n34633 = ~n13318 & n31839;
  assign n34634 = ~n14974 & n34633;
  assign n34635 = n14979 & n34634;
  assign n34636 = ~n34632 & ~n34635;
  assign n34637 = ~n34571 & n34636;
  assign n34638 = ~n13407 & n31835;
  assign n34639 = ~n14467 & n34638;
  assign n34640 = ~n15067 & n34639;
  assign n34641 = n15074 & n34640;
  assign n34642 = ~n13493 & n31900;
  assign n34643 = ~n14467 & n34642;
  assign n34644 = ~n14573 & n34643;
  assign n34645 = ~n15156 & n34644;
  assign n34646 = n15166 & n34645;
  assign n34647 = ~n34641 & ~n34646;
  assign n34648 = n34637 & n34647;
  assign n34649 = ~n12471 & n29527;
  assign n34650 = ~n14467 & n34649;
  assign n34651 = ~n14466 & n34650;
  assign n34652 = n14574 & n34651;
  assign n34653 = n15599 & n34652;
  assign n34654 = n15595 & n34653;
  assign n34655 = n15593 & n34654;
  assign n34656 = n15615 & n34655;
  assign n34657 = ~n12121 & n31789;
  assign n34658 = ~n14467 & n34657;
  assign n34659 = ~n13726 & n34658;
  assign n34660 = n14737 & n34659;
  assign n34661 = n15417 & n34660;
  assign n34662 = n15407 & n34661;
  assign n34663 = ~n34656 & ~n34662;
  assign n34664 = n34648 & n34663;
  assign n34665 = n34565 & n34664;
  assign n34666 = n34541 & n34665;
  assign n34667 = n14981 & n22055;
  assign n34668 = ~n3066 & n34667;
  assign n34669 = ~n3983 & n34668;
  assign n34670 = ~n4003 & n34669;
  assign n34671 = ~n4024 & n34670;
  assign n34672 = ~n4999 & n34671;
  assign n34673 = ~n5827 & n34672;
  assign n34674 = ~n6893 & n34673;
  assign n34675 = ~n7890 & n34674;
  assign n34676 = ~n9131 & n34675;
  assign n34677 = ~n14797 & n34676;
  assign n34678 = ~n14796 & n34677;
  assign n34679 = ~n10278 & n34678;
  assign n34680 = ~n11662 & n34679;
  assign n34681 = ~n14795 & n34680;
  assign n34682 = ~n14794 & n34681;
  assign n34683 = n14817 & n34682;
  assign n34684 = n14820 & n34683;
  assign n34685 = n14824 & n34684;
  assign n34686 = n14793 & n34685;
  assign n34687 = n14847 & n34686;
  assign n34688 = n15386 & n27238;
  assign n34689 = ~n6784 & n34688;
  assign n34690 = ~n7158 & n34689;
  assign n34691 = ~n8250 & n34690;
  assign n34692 = ~n9414 & n34691;
  assign n34693 = ~n15287 & n34692;
  assign n34694 = ~n15286 & n34693;
  assign n34695 = ~n10667 & n34694;
  assign n34696 = ~n12083 & n34695;
  assign n34697 = ~n14467 & n34696;
  assign n34698 = ~n14466 & n34697;
  assign n34699 = n14574 & n34698;
  assign n34700 = n15302 & n34699;
  assign n34701 = n15306 & n34700;
  assign n34702 = n15285 & n34701;
  assign n34703 = n15329 & n34702;
  assign n34704 = pi185 & ~n9913;
  assign n34705 = n15548 & n34704;
  assign n34706 = ~n9929 & n34705;
  assign n34707 = ~n15497 & n34706;
  assign n34708 = ~n15496 & n34707;
  assign n34709 = ~n11266 & n34708;
  assign n34710 = ~n11588 & n34709;
  assign n34711 = ~n14467 & n34710;
  assign n34712 = ~n14466 & n34711;
  assign n34713 = n14574 & n34712;
  assign n34714 = n15508 & n34713;
  assign n34715 = n15512 & n34714;
  assign n34716 = n15495 & n34715;
  assign n34717 = n15535 & n34716;
  assign n34718 = ~n34703 & ~n34717;
  assign n34719 = ~n34687 & n34718;
  assign n34720 = pi105 & ~n4401;
  assign n34721 = n13494 & n34720;
  assign n34722 = ~n4817 & n34721;
  assign n34723 = ~n4902 & n34722;
  assign n34724 = ~n6001 & n34723;
  assign n34725 = ~n7014 & n34724;
  assign n34726 = ~n8114 & n34725;
  assign n34727 = ~n9276 & n34726;
  assign n34728 = ~n15107 & n34727;
  assign n34729 = ~n15106 & n34728;
  assign n34730 = ~n10523 & n34729;
  assign n34731 = ~n11928 & n34730;
  assign n34732 = ~n14467 & n34731;
  assign n34733 = ~n14573 & n34732;
  assign n34734 = n15122 & n34733;
  assign n34735 = n15125 & n34734;
  assign n34736 = n15129 & n34735;
  assign n34737 = n15105 & n34736;
  assign n34738 = n15152 & n34737;
  assign n34739 = pi233 & ~n14416;
  assign n34740 = n15890 & n34739;
  assign n34741 = ~n14519 & n34740;
  assign n34742 = ~n15742 & n34741;
  assign n34743 = ~n14467 & n34742;
  assign n34744 = ~n14466 & n34743;
  assign n34745 = n14574 & n34744;
  assign n34746 = ~n14577 & n34745;
  assign n34747 = n15756 & n34746;
  assign n34748 = n14457 & n34747;
  assign n34749 = n15854 & n34748;
  assign n34750 = ~n34738 & ~n34749;
  assign n34751 = n13408 & n27270;
  assign n34752 = ~n3940 & n34751;
  assign n34753 = ~n4001 & n34752;
  assign n34754 = ~n5043 & n34753;
  assign n34755 = ~n5943 & n34754;
  assign n34756 = ~n6951 & n34755;
  assign n34757 = ~n8037 & n34756;
  assign n34758 = ~n9200 & n34757;
  assign n34759 = ~n15012 & n34758;
  assign n34760 = ~n15011 & n34759;
  assign n34761 = ~n10445 & n34760;
  assign n34762 = ~n11846 & n34761;
  assign n34763 = ~n14467 & n34762;
  assign n34764 = ~n15010 & n34763;
  assign n34765 = n15030 & n34764;
  assign n34766 = n15033 & n34765;
  assign n34767 = n15037 & n34766;
  assign n34768 = n15009 & n34767;
  assign n34769 = n15060 & n34768;
  assign n34770 = pi241 & ~n14568;
  assign n34771 = ~n14520 & n34770;
  assign n34772 = ~n14467 & n34771;
  assign n34773 = ~n14466 & n34772;
  assign n34774 = n14574 & n34773;
  assign n34775 = ~n14465 & n34774;
  assign n34776 = n14581 & n34775;
  assign n34777 = n14457 & n34776;
  assign n34778 = n14715 & n34777;
  assign n34779 = ~n34769 & ~n34778;
  assign n34780 = n34750 & n34779;
  assign n34781 = n15247 & n31984;
  assign n34782 = ~n5808 & n34781;
  assign n34783 = ~n6056 & n34782;
  assign n34784 = ~n7073 & n34783;
  assign n34785 = ~n8179 & n34784;
  assign n34786 = ~n9344 & n34785;
  assign n34787 = ~n15195 & n34786;
  assign n34788 = ~n15194 & n34787;
  assign n34789 = ~n10594 & n34788;
  assign n34790 = ~n12005 & n34789;
  assign n34791 = ~n14467 & n34790;
  assign n34792 = ~n14572 & n34791;
  assign n34793 = n15208 & n34792;
  assign n34794 = n15211 & n34793;
  assign n34795 = n15215 & n34794;
  assign n34796 = n15193 & n34795;
  assign n34797 = n15238 & n34796;
  assign n34798 = n15424 & n23526;
  assign n34799 = ~n7869 & n34798;
  assign n34800 = ~n8346 & n34799;
  assign n34801 = ~n9485 & n34800;
  assign n34802 = ~n15345 & n34801;
  assign n34803 = ~n15344 & n34802;
  assign n34804 = ~n10741 & n34803;
  assign n34805 = ~n12158 & n34804;
  assign n34806 = ~n14467 & n34805;
  assign n34807 = ~n14466 & n34806;
  assign n34808 = n14574 & n34807;
  assign n34809 = n15357 & n34808;
  assign n34810 = n15361 & n34809;
  assign n34811 = n15343 & n34810;
  assign n34812 = n15384 & n34811;
  assign n34813 = ~n34797 & ~n34812;
  assign n34814 = n14858 & n27215;
  assign n34815 = ~n1372 & n34814;
  assign n34816 = ~n2243 & n34815;
  assign n34817 = ~n3104 & n34816;
  assign n34818 = ~n3971 & n34817;
  assign n34819 = ~n4003 & n34818;
  assign n34820 = ~n4872 & n34819;
  assign n34821 = ~n5801 & n34820;
  assign n34822 = ~n6739 & n34821;
  assign n34823 = ~n7807 & n34822;
  assign n34824 = ~n8989 & n34823;
  assign n34825 = ~n10273 & n34824;
  assign n34826 = ~n14857 & n34825;
  assign n34827 = ~n14856 & n34826;
  assign n34828 = ~n11499 & n34827;
  assign n34829 = ~n13076 & n34828;
  assign n34830 = ~n14855 & n34829;
  assign n34831 = ~n14854 & n34830;
  assign n34832 = n14879 & n34831;
  assign n34833 = n14882 & n34832;
  assign n34834 = n14886 & n34833;
  assign n34835 = n14853 & n34834;
  assign n34836 = n14909 & n34835;
  assign n34837 = pi201 & ~n11168;
  assign n34838 = n15698 & n34837;
  assign n34839 = ~n11188 & n34838;
  assign n34840 = ~n15620 & n34839;
  assign n34841 = ~n15619 & n34840;
  assign n34842 = ~n12380 & n34841;
  assign n34843 = ~n14467 & n34842;
  assign n34844 = ~n14466 & n34843;
  assign n34845 = n14574 & n34844;
  assign n34846 = n15629 & n34845;
  assign n34847 = n15633 & n34846;
  assign n34848 = n15595 & n34847;
  assign n34849 = n15656 & n34848;
  assign n34850 = ~n34836 & ~n34849;
  assign n34851 = n34813 & n34850;
  assign n34852 = n34780 & n34851;
  assign n34853 = n34719 & n34852;
  assign po130 = ~n34666 | ~n34853;
  assign n34855 = n13408 & n27506;
  assign n34856 = ~n3940 & n34855;
  assign n34857 = ~n4001 & n34856;
  assign n34858 = ~n5043 & n34857;
  assign n34859 = ~n5943 & n34858;
  assign n34860 = ~n6951 & n34859;
  assign n34861 = ~n8037 & n34860;
  assign n34862 = ~n9200 & n34861;
  assign n34863 = ~n15012 & n34862;
  assign n34864 = ~n15011 & n34863;
  assign n34865 = ~n10445 & n34864;
  assign n34866 = ~n11846 & n34865;
  assign n34867 = ~n14467 & n34866;
  assign n34868 = ~n15010 & n34867;
  assign n34869 = n15030 & n34868;
  assign n34870 = n15033 & n34869;
  assign n34871 = n15037 & n34870;
  assign n34872 = n15009 & n34871;
  assign n34873 = n15060 & n34872;
  assign n34874 = n15247 & n32306;
  assign n34875 = ~n5808 & n34874;
  assign n34876 = ~n6056 & n34875;
  assign n34877 = ~n7073 & n34876;
  assign n34878 = ~n8179 & n34877;
  assign n34879 = ~n9344 & n34878;
  assign n34880 = ~n15195 & n34879;
  assign n34881 = ~n15194 & n34880;
  assign n34882 = ~n10594 & n34881;
  assign n34883 = ~n12005 & n34882;
  assign n34884 = ~n14467 & n34883;
  assign n34885 = ~n14572 & n34884;
  assign n34886 = n15208 & n34885;
  assign n34887 = n15211 & n34886;
  assign n34888 = n15215 & n34887;
  assign n34889 = n15193 & n34888;
  assign n34890 = n15238 & n34889;
  assign n34891 = ~n34873 & ~n34890;
  assign n34892 = ~n14467 & n32388;
  assign n34893 = ~n14466 & n34892;
  assign n34894 = n14574 & n34893;
  assign n34895 = n15859 & n34894;
  assign n34896 = n15862 & n34895;
  assign n34897 = n15595 & n34896;
  assign n34898 = n15885 & n34897;
  assign n34899 = n14749 & n32413;
  assign n34900 = ~n8834 & n34899;
  assign n34901 = ~n10002 & n34900;
  assign n34902 = ~n14747 & n34901;
  assign n34903 = ~n14746 & n34902;
  assign n34904 = ~n11297 & n34903;
  assign n34905 = ~n12240 & n34904;
  assign n34906 = ~n14467 & n34905;
  assign n34907 = ~n14466 & n34906;
  assign n34908 = n14574 & n34907;
  assign n34909 = n14760 & n34908;
  assign n34910 = n14764 & n34909;
  assign n34911 = n14745 & n34910;
  assign n34912 = n14787 & n34911;
  assign n34913 = ~n34898 & ~n34912;
  assign n34914 = n34891 & n34913;
  assign n34915 = ~n11611 & n32107;
  assign n34916 = ~n14467 & n34915;
  assign n34917 = ~n13820 & n34916;
  assign n34918 = ~n14454 & n34917;
  assign n34919 = ~n14455 & n34918;
  assign n34920 = n14738 & n34919;
  assign n34921 = n14730 & n34920;
  assign n34922 = n14723 & n34921;
  assign n34923 = ~n11551 & n32129;
  assign n34924 = ~n14467 & n34923;
  assign n34925 = ~n13906 & n34924;
  assign n34926 = ~n14452 & n34925;
  assign n34927 = n14456 & n34926;
  assign n34928 = n15571 & n34927;
  assign n34929 = n15585 & n34928;
  assign n34930 = ~n12471 & n29864;
  assign n34931 = ~n14467 & n34930;
  assign n34932 = ~n14466 & n34931;
  assign n34933 = n14574 & n34932;
  assign n34934 = n15599 & n34933;
  assign n34935 = n15595 & n34934;
  assign n34936 = n15593 & n34935;
  assign n34937 = n15615 & n34936;
  assign n34938 = ~n34929 & ~n34937;
  assign n34939 = ~n34922 & n34938;
  assign n34940 = ~n13579 & n32221;
  assign n34941 = ~n14467 & n34940;
  assign n34942 = n14574 & n34941;
  assign n34943 = ~n15270 & n34942;
  assign n34944 = n15276 & n34943;
  assign n34945 = n15269 & n34944;
  assign n34946 = pi250 & ~n501;
  assign n34947 = n12872 & n34946;
  assign n34948 = n15973 & n34947;
  assign n34949 = n16069 & n34948;
  assign n34950 = n16063 & n34949;
  assign n34951 = n16088 & n34950;
  assign n34952 = ~n1172 & n34951;
  assign n34953 = ~n996 & n34952;
  assign n34954 = ~n2306 & n34953;
  assign n34955 = ~n500 & n34954;
  assign n34956 = n16094 & n34955;
  assign n34957 = n16016 & n34956;
  assign n34958 = n16054 & n34957;
  assign n34959 = n16113 & n34958;
  assign n34960 = n16184 & n34959;
  assign n34961 = n16048 & n34960;
  assign n34962 = ~n7236 & n34961;
  assign n34963 = ~n6137 & n34962;
  assign n34964 = n6193 & n34963;
  assign n34965 = n6134 & n34964;
  assign n34966 = ~n8867 & n34965;
  assign n34967 = ~n7235 & n34966;
  assign n34968 = n7296 & n34967;
  assign n34969 = n7231 & n34968;
  assign n34970 = ~n10027 & n34969;
  assign n34971 = ~n8866 & n34970;
  assign n34972 = n8898 & n34971;
  assign n34973 = n8863 & n34972;
  assign n34974 = pi258 & ~n501;
  assign n34975 = n12872 & n34974;
  assign n34976 = n15973 & n34975;
  assign n34977 = n15980 & n34976;
  assign n34978 = n15972 & n34977;
  assign n34979 = n16005 & n34978;
  assign n34980 = ~n1172 & n34979;
  assign n34981 = ~n996 & n34980;
  assign n34982 = ~n2306 & n34981;
  assign n34983 = ~n500 & n34982;
  assign n34984 = n16011 & n34983;
  assign n34985 = n16014 & n34984;
  assign n34986 = n16017 & n34985;
  assign n34987 = n16038 & n34986;
  assign n34988 = n15963 & n34987;
  assign n34989 = n15954 & n34988;
  assign n34990 = ~n7236 & n34989;
  assign n34991 = ~n6137 & n34990;
  assign n34992 = n6193 & n34991;
  assign n34993 = n6134 & n34992;
  assign n34994 = ~n8867 & n34993;
  assign n34995 = ~n7235 & n34994;
  assign n34996 = n7296 & n34995;
  assign n34997 = n7231 & n34996;
  assign n34998 = ~n10027 & n34997;
  assign n34999 = ~n8866 & n34998;
  assign n35000 = n8898 & n34999;
  assign n35001 = n8863 & n35000;
  assign n35002 = ~n34973 & ~n35001;
  assign n35003 = ~n10788 & ~n35002;
  assign n35004 = ~n10026 & n35003;
  assign n35005 = n10072 & n35004;
  assign n35006 = n10021 & n35005;
  assign n35007 = ~n13318 & n32155;
  assign n35008 = ~n14974 & n35007;
  assign n35009 = n14979 & n35008;
  assign n35010 = ~n35006 & ~n35009;
  assign n35011 = ~n34945 & n35010;
  assign n35012 = ~n13407 & n32151;
  assign n35013 = ~n14467 & n35012;
  assign n35014 = ~n15067 & n35013;
  assign n35015 = n15074 & n35014;
  assign n35016 = ~n13493 & n32216;
  assign n35017 = ~n14467 & n35016;
  assign n35018 = ~n14573 & n35017;
  assign n35019 = ~n15156 & n35018;
  assign n35020 = n15166 & n35019;
  assign n35021 = ~n35015 & ~n35020;
  assign n35022 = n35011 & n35021;
  assign n35023 = ~n12181 & n32122;
  assign n35024 = ~n14467 & n35023;
  assign n35025 = ~n13764 & n35024;
  assign n35026 = ~n14455 & n35025;
  assign n35027 = n14737 & n35026;
  assign n35028 = n15463 & n35027;
  assign n35029 = n15452 & n35028;
  assign n35030 = ~n12121 & n32114;
  assign n35031 = ~n14467 & n35030;
  assign n35032 = ~n13726 & n35031;
  assign n35033 = n14737 & n35032;
  assign n35034 = n15417 & n35033;
  assign n35035 = n15407 & n35034;
  assign n35036 = ~n35029 & ~n35035;
  assign n35037 = n35022 & n35036;
  assign n35038 = n34939 & n35037;
  assign n35039 = n34914 & n35038;
  assign n35040 = n14981 & n22280;
  assign n35041 = ~n3066 & n35040;
  assign n35042 = ~n3983 & n35041;
  assign n35043 = ~n4003 & n35042;
  assign n35044 = ~n4024 & n35043;
  assign n35045 = ~n4999 & n35044;
  assign n35046 = ~n5827 & n35045;
  assign n35047 = ~n6893 & n35046;
  assign n35048 = ~n7890 & n35047;
  assign n35049 = ~n9131 & n35048;
  assign n35050 = ~n14797 & n35049;
  assign n35051 = ~n14796 & n35050;
  assign n35052 = ~n10278 & n35051;
  assign n35053 = ~n11662 & n35052;
  assign n35054 = ~n14795 & n35053;
  assign n35055 = ~n14794 & n35054;
  assign n35056 = n14817 & n35055;
  assign n35057 = n14820 & n35056;
  assign n35058 = n14824 & n35057;
  assign n35059 = n14793 & n35058;
  assign n35060 = n14847 & n35059;
  assign n35061 = n15386 & n27435;
  assign n35062 = ~n6784 & n35061;
  assign n35063 = ~n7158 & n35062;
  assign n35064 = ~n8250 & n35063;
  assign n35065 = ~n9414 & n35064;
  assign n35066 = ~n15287 & n35065;
  assign n35067 = ~n15286 & n35066;
  assign n35068 = ~n10667 & n35067;
  assign n35069 = ~n12083 & n35068;
  assign n35070 = ~n14467 & n35069;
  assign n35071 = ~n14466 & n35070;
  assign n35072 = n14574 & n35071;
  assign n35073 = n15302 & n35072;
  assign n35074 = n15306 & n35073;
  assign n35075 = n15285 & n35074;
  assign n35076 = n15329 & n35075;
  assign n35077 = pi186 & ~n9913;
  assign n35078 = n15548 & n35077;
  assign n35079 = ~n9929 & n35078;
  assign n35080 = ~n15497 & n35079;
  assign n35081 = ~n15496 & n35080;
  assign n35082 = ~n11266 & n35081;
  assign n35083 = ~n11588 & n35082;
  assign n35084 = ~n14467 & n35083;
  assign n35085 = ~n14466 & n35084;
  assign n35086 = n14574 & n35085;
  assign n35087 = n15508 & n35086;
  assign n35088 = n15512 & n35087;
  assign n35089 = n15495 & n35088;
  assign n35090 = n15535 & n35089;
  assign n35091 = ~n35076 & ~n35090;
  assign n35092 = ~n35060 & n35091;
  assign n35093 = pi234 & ~n14416;
  assign n35094 = n15890 & n35093;
  assign n35095 = ~n14519 & n35094;
  assign n35096 = ~n15742 & n35095;
  assign n35097 = ~n14467 & n35096;
  assign n35098 = ~n14466 & n35097;
  assign n35099 = n14574 & n35098;
  assign n35100 = ~n14577 & n35099;
  assign n35101 = n15756 & n35100;
  assign n35102 = n14457 & n35101;
  assign n35103 = n15854 & n35102;
  assign n35104 = n14858 & n27477;
  assign n35105 = ~n1372 & n35104;
  assign n35106 = ~n2243 & n35105;
  assign n35107 = ~n3104 & n35106;
  assign n35108 = ~n3971 & n35107;
  assign n35109 = ~n4003 & n35108;
  assign n35110 = ~n4872 & n35109;
  assign n35111 = ~n5801 & n35110;
  assign n35112 = ~n6739 & n35111;
  assign n35113 = ~n7807 & n35112;
  assign n35114 = ~n8989 & n35113;
  assign n35115 = ~n10273 & n35114;
  assign n35116 = ~n14857 & n35115;
  assign n35117 = ~n14856 & n35116;
  assign n35118 = ~n11499 & n35117;
  assign n35119 = ~n13076 & n35118;
  assign n35120 = ~n14855 & n35119;
  assign n35121 = ~n14854 & n35120;
  assign n35122 = n14879 & n35121;
  assign n35123 = n14882 & n35122;
  assign n35124 = n14886 & n35123;
  assign n35125 = n14853 & n35124;
  assign n35126 = n14909 & n35125;
  assign n35127 = ~n35103 & ~n35126;
  assign n35128 = pi106 & ~n4401;
  assign n35129 = n13494 & n35128;
  assign n35130 = ~n4817 & n35129;
  assign n35131 = ~n4902 & n35130;
  assign n35132 = ~n6001 & n35131;
  assign n35133 = ~n7014 & n35132;
  assign n35134 = ~n8114 & n35133;
  assign n35135 = ~n9276 & n35134;
  assign n35136 = ~n15107 & n35135;
  assign n35137 = ~n15106 & n35136;
  assign n35138 = ~n10523 & n35137;
  assign n35139 = ~n11928 & n35138;
  assign n35140 = ~n14467 & n35139;
  assign n35141 = ~n14573 & n35140;
  assign n35142 = n15122 & n35141;
  assign n35143 = n15125 & n35142;
  assign n35144 = n15129 & n35143;
  assign n35145 = n15105 & n35144;
  assign n35146 = n15152 & n35145;
  assign n35147 = pi058 & ~n1740;
  assign n35148 = n13259 & n35147;
  assign n35149 = ~n2242 & n35148;
  assign n35150 = ~n3095 & n35149;
  assign n35151 = ~n3997 & n35150;
  assign n35152 = ~n4003 & n35151;
  assign n35153 = ~n4837 & n35152;
  assign n35154 = ~n5822 & n35153;
  assign n35155 = ~n6820 & n35154;
  assign n35156 = ~n7785 & n35155;
  assign n35157 = ~n9027 & n35156;
  assign n35158 = ~n10245 & n35157;
  assign n35159 = ~n14919 & n35158;
  assign n35160 = ~n14918 & n35159;
  assign n35161 = ~n11536 & n35160;
  assign n35162 = ~n13036 & n35161;
  assign n35163 = ~n14917 & n35162;
  assign n35164 = ~n14916 & n35163;
  assign n35165 = n14940 & n35164;
  assign n35166 = n14943 & n35165;
  assign n35167 = n14947 & n35166;
  assign n35168 = n14915 & n35167;
  assign n35169 = n14970 & n35168;
  assign n35170 = ~n35146 & ~n35169;
  assign n35171 = n35127 & n35170;
  assign n35172 = pi242 & ~n14568;
  assign n35173 = ~n14520 & n35172;
  assign n35174 = ~n14467 & n35173;
  assign n35175 = ~n14466 & n35174;
  assign n35176 = n14574 & n35175;
  assign n35177 = ~n14465 & n35176;
  assign n35178 = n14581 & n35177;
  assign n35179 = n14457 & n35178;
  assign n35180 = n14715 & n35179;
  assign n35181 = n15424 & n23752;
  assign n35182 = ~n7869 & n35181;
  assign n35183 = ~n8346 & n35182;
  assign n35184 = ~n9485 & n35183;
  assign n35185 = ~n15345 & n35184;
  assign n35186 = ~n15344 & n35185;
  assign n35187 = ~n10741 & n35186;
  assign n35188 = ~n12158 & n35187;
  assign n35189 = ~n14467 & n35188;
  assign n35190 = ~n14466 & n35189;
  assign n35191 = n14574 & n35190;
  assign n35192 = n15357 & n35191;
  assign n35193 = n15361 & n35192;
  assign n35194 = n15343 & n35193;
  assign n35195 = n15384 & n35194;
  assign n35196 = ~n35180 & ~n35195;
  assign n35197 = pi202 & ~n11168;
  assign n35198 = n15698 & n35197;
  assign n35199 = ~n11188 & n35198;
  assign n35200 = ~n15620 & n35199;
  assign n35201 = ~n15619 & n35200;
  assign n35202 = ~n12380 & n35201;
  assign n35203 = ~n14467 & n35202;
  assign n35204 = ~n14466 & n35203;
  assign n35205 = n14574 & n35204;
  assign n35206 = n15629 & n35205;
  assign n35207 = n15633 & n35206;
  assign n35208 = n15595 & n35207;
  assign n35209 = n15656 & n35208;
  assign n35210 = pi218 & ~n12841;
  assign n35211 = n12775 & n35210;
  assign n35212 = ~n12902 & n35211;
  assign n35213 = ~n15659 & n35212;
  assign n35214 = ~n15658 & n35213;
  assign n35215 = ~n14467 & n35214;
  assign n35216 = ~n14466 & n35215;
  assign n35217 = n14574 & n35216;
  assign n35218 = n15666 & n35217;
  assign n35219 = n15669 & n35218;
  assign n35220 = n15595 & n35219;
  assign n35221 = n15692 & n35220;
  assign n35222 = ~n35209 & ~n35221;
  assign n35223 = n35196 & n35222;
  assign n35224 = n35171 & n35223;
  assign n35225 = n35092 & n35224;
  assign po131 = ~n35039 | ~n35225;
  assign n35227 = n14858 & n27731;
  assign n35228 = ~n1372 & n35227;
  assign n35229 = ~n2243 & n35228;
  assign n35230 = ~n3104 & n35229;
  assign n35231 = ~n3971 & n35230;
  assign n35232 = ~n4003 & n35231;
  assign n35233 = ~n4872 & n35232;
  assign n35234 = ~n5801 & n35233;
  assign n35235 = ~n6739 & n35234;
  assign n35236 = ~n7807 & n35235;
  assign n35237 = ~n8989 & n35236;
  assign n35238 = ~n10273 & n35237;
  assign n35239 = ~n14857 & n35238;
  assign n35240 = ~n14856 & n35239;
  assign n35241 = ~n11499 & n35240;
  assign n35242 = ~n13076 & n35241;
  assign n35243 = ~n14855 & n35242;
  assign n35244 = ~n14854 & n35243;
  assign n35245 = n14879 & n35244;
  assign n35246 = n14882 & n35245;
  assign n35247 = n14886 & n35246;
  assign n35248 = n14853 & n35247;
  assign n35249 = n14909 & n35248;
  assign n35250 = ~n14467 & n32576;
  assign n35251 = ~n14466 & n35250;
  assign n35252 = n14574 & n35251;
  assign n35253 = n15859 & n35252;
  assign n35254 = n15862 & n35253;
  assign n35255 = n15595 & n35254;
  assign n35256 = n15885 & n35255;
  assign n35257 = ~n35249 & ~n35256;
  assign n35258 = n15424 & n23945;
  assign n35259 = ~n7869 & n35258;
  assign n35260 = ~n8346 & n35259;
  assign n35261 = ~n9485 & n35260;
  assign n35262 = ~n15345 & n35261;
  assign n35263 = ~n15344 & n35262;
  assign n35264 = ~n10741 & n35263;
  assign n35265 = ~n12158 & n35264;
  assign n35266 = ~n14467 & n35265;
  assign n35267 = ~n14466 & n35266;
  assign n35268 = n14574 & n35267;
  assign n35269 = n15357 & n35268;
  assign n35270 = n15361 & n35269;
  assign n35271 = n15343 & n35270;
  assign n35272 = n15384 & n35271;
  assign n35273 = n15247 & n32586;
  assign n35274 = ~n5808 & n35273;
  assign n35275 = ~n6056 & n35274;
  assign n35276 = ~n7073 & n35275;
  assign n35277 = ~n8179 & n35276;
  assign n35278 = ~n9344 & n35277;
  assign n35279 = ~n15195 & n35278;
  assign n35280 = ~n15194 & n35279;
  assign n35281 = ~n10594 & n35280;
  assign n35282 = ~n12005 & n35281;
  assign n35283 = ~n14467 & n35282;
  assign n35284 = ~n14572 & n35283;
  assign n35285 = n15208 & n35284;
  assign n35286 = n15211 & n35285;
  assign n35287 = n15215 & n35286;
  assign n35288 = n15193 & n35287;
  assign n35289 = n15238 & n35288;
  assign n35290 = ~n35272 & ~n35289;
  assign n35291 = n35257 & n35290;
  assign n35292 = ~n12181 & n32447;
  assign n35293 = ~n14467 & n35292;
  assign n35294 = ~n13764 & n35293;
  assign n35295 = ~n14455 & n35294;
  assign n35296 = n14737 & n35295;
  assign n35297 = n15463 & n35296;
  assign n35298 = n15452 & n35297;
  assign n35299 = ~n11611 & n32454;
  assign n35300 = ~n14467 & n35299;
  assign n35301 = ~n13820 & n35300;
  assign n35302 = ~n14454 & n35301;
  assign n35303 = ~n14455 & n35302;
  assign n35304 = n14738 & n35303;
  assign n35305 = n14730 & n35304;
  assign n35306 = n14723 & n35305;
  assign n35307 = ~n11551 & n32432;
  assign n35308 = ~n14467 & n35307;
  assign n35309 = ~n13906 & n35308;
  assign n35310 = ~n14452 & n35309;
  assign n35311 = n14456 & n35310;
  assign n35312 = n15571 & n35311;
  assign n35313 = n15585 & n35312;
  assign n35314 = ~n35306 & ~n35313;
  assign n35315 = ~n35298 & n35314;
  assign n35316 = ~n13407 & n32485;
  assign n35317 = ~n14467 & n35316;
  assign n35318 = ~n15067 & n35317;
  assign n35319 = n15074 & n35318;
  assign n35320 = ~n13318 & n32489;
  assign n35321 = ~n14974 & n35320;
  assign n35322 = n14979 & n35321;
  assign n35323 = pi259 & ~n501;
  assign n35324 = n12872 & n35323;
  assign n35325 = n15973 & n35324;
  assign n35326 = n15980 & n35325;
  assign n35327 = n15972 & n35326;
  assign n35328 = n16005 & n35327;
  assign n35329 = ~n1172 & n35328;
  assign n35330 = ~n996 & n35329;
  assign n35331 = ~n2306 & n35330;
  assign n35332 = ~n500 & n35331;
  assign n35333 = n16011 & n35332;
  assign n35334 = n16014 & n35333;
  assign n35335 = n16017 & n35334;
  assign n35336 = n16038 & n35335;
  assign n35337 = n15963 & n35336;
  assign n35338 = n15954 & n35337;
  assign n35339 = ~n7236 & n35338;
  assign n35340 = ~n6137 & n35339;
  assign n35341 = n6193 & n35340;
  assign n35342 = n6134 & n35341;
  assign n35343 = ~n8867 & n35342;
  assign n35344 = ~n7235 & n35343;
  assign n35345 = n7296 & n35344;
  assign n35346 = n7231 & n35345;
  assign n35347 = ~n10027 & n35346;
  assign n35348 = ~n8866 & n35347;
  assign n35349 = n8898 & n35348;
  assign n35350 = n8863 & n35349;
  assign n35351 = pi251 & ~n501;
  assign n35352 = n12872 & n35351;
  assign n35353 = n15973 & n35352;
  assign n35354 = n16069 & n35353;
  assign n35355 = n16063 & n35354;
  assign n35356 = n16088 & n35355;
  assign n35357 = ~n1172 & n35356;
  assign n35358 = ~n996 & n35357;
  assign n35359 = ~n2306 & n35358;
  assign n35360 = ~n500 & n35359;
  assign n35361 = n16094 & n35360;
  assign n35362 = n16016 & n35361;
  assign n35363 = n16054 & n35362;
  assign n35364 = n16113 & n35363;
  assign n35365 = n16184 & n35364;
  assign n35366 = n16048 & n35365;
  assign n35367 = ~n7236 & n35366;
  assign n35368 = ~n6137 & n35367;
  assign n35369 = n6193 & n35368;
  assign n35370 = n6134 & n35369;
  assign n35371 = ~n8867 & n35370;
  assign n35372 = ~n7235 & n35371;
  assign n35373 = n7296 & n35372;
  assign n35374 = n7231 & n35373;
  assign n35375 = ~n10027 & n35374;
  assign n35376 = ~n8866 & n35375;
  assign n35377 = n8898 & n35376;
  assign n35378 = n8863 & n35377;
  assign n35379 = ~n35350 & ~n35378;
  assign n35380 = ~n10788 & ~n35379;
  assign n35381 = ~n10026 & n35380;
  assign n35382 = n10072 & n35381;
  assign n35383 = n10021 & n35382;
  assign n35384 = ~n35322 & ~n35383;
  assign n35385 = ~n35319 & n35384;
  assign n35386 = ~n13493 & n32550;
  assign n35387 = ~n14467 & n35386;
  assign n35388 = ~n14573 & n35387;
  assign n35389 = ~n15156 & n35388;
  assign n35390 = n15166 & n35389;
  assign n35391 = ~n13579 & n32555;
  assign n35392 = ~n14467 & n35391;
  assign n35393 = n14574 & n35392;
  assign n35394 = ~n15270 & n35393;
  assign n35395 = n15276 & n35394;
  assign n35396 = n15269 & n35395;
  assign n35397 = ~n35390 & ~n35396;
  assign n35398 = n35385 & n35397;
  assign n35399 = ~n12471 & n30085;
  assign n35400 = ~n14467 & n35399;
  assign n35401 = ~n14466 & n35400;
  assign n35402 = n14574 & n35401;
  assign n35403 = n15599 & n35402;
  assign n35404 = n15595 & n35403;
  assign n35405 = n15593 & n35404;
  assign n35406 = n15615 & n35405;
  assign n35407 = ~n12121 & n32439;
  assign n35408 = ~n14467 & n35407;
  assign n35409 = ~n13726 & n35408;
  assign n35410 = n14737 & n35409;
  assign n35411 = n15417 & n35410;
  assign n35412 = n15407 & n35411;
  assign n35413 = ~n35406 & ~n35412;
  assign n35414 = n35398 & n35413;
  assign n35415 = n35315 & n35414;
  assign n35416 = n35291 & n35415;
  assign n35417 = n14981 & n22447;
  assign n35418 = ~n3066 & n35417;
  assign n35419 = ~n3983 & n35418;
  assign n35420 = ~n4003 & n35419;
  assign n35421 = ~n4024 & n35420;
  assign n35422 = ~n4999 & n35421;
  assign n35423 = ~n5827 & n35422;
  assign n35424 = ~n6893 & n35423;
  assign n35425 = ~n7890 & n35424;
  assign n35426 = ~n9131 & n35425;
  assign n35427 = ~n14797 & n35426;
  assign n35428 = ~n14796 & n35427;
  assign n35429 = ~n10278 & n35428;
  assign n35430 = ~n11662 & n35429;
  assign n35431 = ~n14795 & n35430;
  assign n35432 = ~n14794 & n35431;
  assign n35433 = n14817 & n35432;
  assign n35434 = n14820 & n35433;
  assign n35435 = n14824 & n35434;
  assign n35436 = n14793 & n35435;
  assign n35437 = n14847 & n35436;
  assign n35438 = pi219 & ~n12841;
  assign n35439 = n12775 & n35438;
  assign n35440 = ~n12902 & n35439;
  assign n35441 = ~n15659 & n35440;
  assign n35442 = ~n15658 & n35441;
  assign n35443 = ~n14467 & n35442;
  assign n35444 = ~n14466 & n35443;
  assign n35445 = n14574 & n35444;
  assign n35446 = n15666 & n35445;
  assign n35447 = n15669 & n35446;
  assign n35448 = n15595 & n35447;
  assign n35449 = n15692 & n35448;
  assign n35450 = pi187 & ~n9913;
  assign n35451 = n15548 & n35450;
  assign n35452 = ~n9929 & n35451;
  assign n35453 = ~n15497 & n35452;
  assign n35454 = ~n15496 & n35453;
  assign n35455 = ~n11266 & n35454;
  assign n35456 = ~n11588 & n35455;
  assign n35457 = ~n14467 & n35456;
  assign n35458 = ~n14466 & n35457;
  assign n35459 = n14574 & n35458;
  assign n35460 = n15508 & n35459;
  assign n35461 = n15512 & n35460;
  assign n35462 = n15495 & n35461;
  assign n35463 = n15535 & n35462;
  assign n35464 = ~n35449 & ~n35463;
  assign n35465 = ~n35437 & n35464;
  assign n35466 = n14749 & n32725;
  assign n35467 = ~n8834 & n35466;
  assign n35468 = ~n10002 & n35467;
  assign n35469 = ~n14747 & n35468;
  assign n35470 = ~n14746 & n35469;
  assign n35471 = ~n11297 & n35470;
  assign n35472 = ~n12240 & n35471;
  assign n35473 = ~n14467 & n35472;
  assign n35474 = ~n14466 & n35473;
  assign n35475 = n14574 & n35474;
  assign n35476 = n14760 & n35475;
  assign n35477 = n14764 & n35476;
  assign n35478 = n14745 & n35477;
  assign n35479 = n14787 & n35478;
  assign n35480 = pi107 & ~n4401;
  assign n35481 = n13494 & n35480;
  assign n35482 = ~n4817 & n35481;
  assign n35483 = ~n4902 & n35482;
  assign n35484 = ~n6001 & n35483;
  assign n35485 = ~n7014 & n35484;
  assign n35486 = ~n8114 & n35485;
  assign n35487 = ~n9276 & n35486;
  assign n35488 = ~n15107 & n35487;
  assign n35489 = ~n15106 & n35488;
  assign n35490 = ~n10523 & n35489;
  assign n35491 = ~n11928 & n35490;
  assign n35492 = ~n14467 & n35491;
  assign n35493 = ~n14573 & n35492;
  assign n35494 = n15122 & n35493;
  assign n35495 = n15125 & n35494;
  assign n35496 = n15129 & n35495;
  assign n35497 = n15105 & n35496;
  assign n35498 = n15152 & n35497;
  assign n35499 = ~n35479 & ~n35498;
  assign n35500 = pi243 & ~n14568;
  assign n35501 = ~n14520 & n35500;
  assign n35502 = ~n14467 & n35501;
  assign n35503 = ~n14466 & n35502;
  assign n35504 = n14574 & n35503;
  assign n35505 = ~n14465 & n35504;
  assign n35506 = n14581 & n35505;
  assign n35507 = n14457 & n35506;
  assign n35508 = n14715 & n35507;
  assign n35509 = pi203 & ~n11168;
  assign n35510 = n15698 & n35509;
  assign n35511 = ~n11188 & n35510;
  assign n35512 = ~n15620 & n35511;
  assign n35513 = ~n15619 & n35512;
  assign n35514 = ~n12380 & n35513;
  assign n35515 = ~n14467 & n35514;
  assign n35516 = ~n14466 & n35515;
  assign n35517 = n14574 & n35516;
  assign n35518 = n15629 & n35517;
  assign n35519 = n15633 & n35518;
  assign n35520 = n15595 & n35519;
  assign n35521 = n15656 & n35520;
  assign n35522 = ~n35508 & ~n35521;
  assign n35523 = n35499 & n35522;
  assign n35524 = pi059 & ~n1740;
  assign n35525 = n13259 & n35524;
  assign n35526 = ~n2242 & n35525;
  assign n35527 = ~n3095 & n35526;
  assign n35528 = ~n3997 & n35527;
  assign n35529 = ~n4003 & n35528;
  assign n35530 = ~n4837 & n35529;
  assign n35531 = ~n5822 & n35530;
  assign n35532 = ~n6820 & n35531;
  assign n35533 = ~n7785 & n35532;
  assign n35534 = ~n9027 & n35533;
  assign n35535 = ~n10245 & n35534;
  assign n35536 = ~n14919 & n35535;
  assign n35537 = ~n14918 & n35536;
  assign n35538 = ~n11536 & n35537;
  assign n35539 = ~n13036 & n35538;
  assign n35540 = ~n14917 & n35539;
  assign n35541 = ~n14916 & n35540;
  assign n35542 = n14940 & n35541;
  assign n35543 = n14943 & n35542;
  assign n35544 = n14947 & n35543;
  assign n35545 = n14915 & n35544;
  assign n35546 = n14970 & n35545;
  assign n35547 = n13408 & n27770;
  assign n35548 = ~n3940 & n35547;
  assign n35549 = ~n4001 & n35548;
  assign n35550 = ~n5043 & n35549;
  assign n35551 = ~n5943 & n35550;
  assign n35552 = ~n6951 & n35551;
  assign n35553 = ~n8037 & n35552;
  assign n35554 = ~n9200 & n35553;
  assign n35555 = ~n15012 & n35554;
  assign n35556 = ~n15011 & n35555;
  assign n35557 = ~n10445 & n35556;
  assign n35558 = ~n11846 & n35557;
  assign n35559 = ~n14467 & n35558;
  assign n35560 = ~n15010 & n35559;
  assign n35561 = n15030 & n35560;
  assign n35562 = n15033 & n35561;
  assign n35563 = n15037 & n35562;
  assign n35564 = n15009 & n35563;
  assign n35565 = n15060 & n35564;
  assign n35566 = ~n35546 & ~n35565;
  assign n35567 = n15386 & n27789;
  assign n35568 = ~n6784 & n35567;
  assign n35569 = ~n7158 & n35568;
  assign n35570 = ~n8250 & n35569;
  assign n35571 = ~n9414 & n35570;
  assign n35572 = ~n15287 & n35571;
  assign n35573 = ~n15286 & n35572;
  assign n35574 = ~n10667 & n35573;
  assign n35575 = ~n12083 & n35574;
  assign n35576 = ~n14467 & n35575;
  assign n35577 = ~n14466 & n35576;
  assign n35578 = n14574 & n35577;
  assign n35579 = n15302 & n35578;
  assign n35580 = n15306 & n35579;
  assign n35581 = n15285 & n35580;
  assign n35582 = n15329 & n35581;
  assign n35583 = pi235 & ~n14416;
  assign n35584 = n15890 & n35583;
  assign n35585 = ~n14519 & n35584;
  assign n35586 = ~n15742 & n35585;
  assign n35587 = ~n14467 & n35586;
  assign n35588 = ~n14466 & n35587;
  assign n35589 = n14574 & n35588;
  assign n35590 = ~n14577 & n35589;
  assign n35591 = n15756 & n35590;
  assign n35592 = n14457 & n35591;
  assign n35593 = n15854 & n35592;
  assign n35594 = ~n35582 & ~n35593;
  assign n35595 = n35566 & n35594;
  assign n35596 = n35523 & n35595;
  assign n35597 = n35465 & n35596;
  assign po132 = ~n35416 | ~n35597;
  assign n35599 = pi060 & ~n1740;
  assign n35600 = n13259 & n35599;
  assign n35601 = ~n2242 & n35600;
  assign n35602 = ~n3095 & n35601;
  assign n35603 = ~n3997 & n35602;
  assign n35604 = ~n4003 & n35603;
  assign n35605 = ~n4837 & n35604;
  assign n35606 = ~n5822 & n35605;
  assign n35607 = ~n6820 & n35606;
  assign n35608 = ~n7785 & n35607;
  assign n35609 = ~n9027 & n35608;
  assign n35610 = ~n10245 & n35609;
  assign n35611 = ~n14919 & n35610;
  assign n35612 = ~n14918 & n35611;
  assign n35613 = ~n11536 & n35612;
  assign n35614 = ~n13036 & n35613;
  assign n35615 = ~n14917 & n35614;
  assign n35616 = ~n14916 & n35615;
  assign n35617 = n14940 & n35616;
  assign n35618 = n14943 & n35617;
  assign n35619 = n14947 & n35618;
  assign n35620 = n14915 & n35619;
  assign n35621 = n14970 & n35620;
  assign n35622 = pi244 & ~n14568;
  assign n35623 = ~n14520 & n35622;
  assign n35624 = ~n14467 & n35623;
  assign n35625 = ~n14466 & n35624;
  assign n35626 = n14574 & n35625;
  assign n35627 = ~n14465 & n35626;
  assign n35628 = n14581 & n35627;
  assign n35629 = n14457 & n35628;
  assign n35630 = n14715 & n35629;
  assign n35631 = ~n35621 & ~n35630;
  assign n35632 = pi204 & ~n11168;
  assign n35633 = n15698 & n35632;
  assign n35634 = ~n11188 & n35633;
  assign n35635 = ~n15620 & n35634;
  assign n35636 = ~n15619 & n35635;
  assign n35637 = ~n12380 & n35636;
  assign n35638 = ~n14467 & n35637;
  assign n35639 = ~n14466 & n35638;
  assign n35640 = n14574 & n35639;
  assign n35641 = n15629 & n35640;
  assign n35642 = n15633 & n35641;
  assign n35643 = n15595 & n35642;
  assign n35644 = n15656 & n35643;
  assign n35645 = pi220 & ~n12841;
  assign n35646 = n12775 & n35645;
  assign n35647 = ~n12902 & n35646;
  assign n35648 = ~n15659 & n35647;
  assign n35649 = ~n15658 & n35648;
  assign n35650 = ~n14467 & n35649;
  assign n35651 = ~n14466 & n35650;
  assign n35652 = n14574 & n35651;
  assign n35653 = n15666 & n35652;
  assign n35654 = n15669 & n35653;
  assign n35655 = n15595 & n35654;
  assign n35656 = n15692 & n35655;
  assign n35657 = ~n35644 & ~n35656;
  assign n35658 = n35631 & n35657;
  assign n35659 = ~n11551 & n32779;
  assign n35660 = ~n14467 & n35659;
  assign n35661 = ~n13906 & n35660;
  assign n35662 = ~n14452 & n35661;
  assign n35663 = n14456 & n35662;
  assign n35664 = n15571 & n35663;
  assign n35665 = n15585 & n35664;
  assign n35666 = ~n12181 & n32764;
  assign n35667 = ~n14467 & n35666;
  assign n35668 = ~n13764 & n35667;
  assign n35669 = ~n14455 & n35668;
  assign n35670 = n14737 & n35669;
  assign n35671 = n15463 & n35670;
  assign n35672 = n15452 & n35671;
  assign n35673 = ~n12121 & n32757;
  assign n35674 = ~n14467 & n35673;
  assign n35675 = ~n13726 & n35674;
  assign n35676 = n14737 & n35675;
  assign n35677 = n15417 & n35676;
  assign n35678 = n15407 & n35677;
  assign n35679 = ~n35672 & ~n35678;
  assign n35680 = ~n35665 & n35679;
  assign n35681 = ~n13407 & n32801;
  assign n35682 = ~n14467 & n35681;
  assign n35683 = ~n15067 & n35682;
  assign n35684 = n15074 & n35683;
  assign n35685 = ~n13318 & n32805;
  assign n35686 = ~n14974 & n35685;
  assign n35687 = n14979 & n35686;
  assign n35688 = pi252 & ~n501;
  assign n35689 = n12872 & n35688;
  assign n35690 = n15973 & n35689;
  assign n35691 = n16069 & n35690;
  assign n35692 = n16063 & n35691;
  assign n35693 = n16088 & n35692;
  assign n35694 = ~n1172 & n35693;
  assign n35695 = ~n996 & n35694;
  assign n35696 = ~n2306 & n35695;
  assign n35697 = ~n500 & n35696;
  assign n35698 = n16094 & n35697;
  assign n35699 = n16016 & n35698;
  assign n35700 = n16054 & n35699;
  assign n35701 = n16113 & n35700;
  assign n35702 = n16184 & n35701;
  assign n35703 = n16048 & n35702;
  assign n35704 = ~n7236 & n35703;
  assign n35705 = ~n6137 & n35704;
  assign n35706 = n6193 & n35705;
  assign n35707 = n6134 & n35706;
  assign n35708 = ~n8867 & n35707;
  assign n35709 = ~n7235 & n35708;
  assign n35710 = n7296 & n35709;
  assign n35711 = n7231 & n35710;
  assign n35712 = ~n10027 & n35711;
  assign n35713 = ~n8866 & n35712;
  assign n35714 = n8898 & n35713;
  assign n35715 = n8863 & n35714;
  assign n35716 = pi260 & ~n501;
  assign n35717 = n12872 & n35716;
  assign n35718 = n15973 & n35717;
  assign n35719 = n15980 & n35718;
  assign n35720 = n15972 & n35719;
  assign n35721 = n16005 & n35720;
  assign n35722 = ~n1172 & n35721;
  assign n35723 = ~n996 & n35722;
  assign n35724 = ~n2306 & n35723;
  assign n35725 = ~n500 & n35724;
  assign n35726 = n16011 & n35725;
  assign n35727 = n16014 & n35726;
  assign n35728 = n16017 & n35727;
  assign n35729 = n16038 & n35728;
  assign n35730 = n15963 & n35729;
  assign n35731 = n15954 & n35730;
  assign n35732 = ~n7236 & n35731;
  assign n35733 = ~n6137 & n35732;
  assign n35734 = n6193 & n35733;
  assign n35735 = n6134 & n35734;
  assign n35736 = ~n8867 & n35735;
  assign n35737 = ~n7235 & n35736;
  assign n35738 = n7296 & n35737;
  assign n35739 = n7231 & n35738;
  assign n35740 = ~n10027 & n35739;
  assign n35741 = ~n8866 & n35740;
  assign n35742 = n8898 & n35741;
  assign n35743 = n8863 & n35742;
  assign n35744 = ~n35715 & ~n35743;
  assign n35745 = ~n10788 & ~n35744;
  assign n35746 = ~n10026 & n35745;
  assign n35747 = n10072 & n35746;
  assign n35748 = n10021 & n35747;
  assign n35749 = ~n35687 & ~n35748;
  assign n35750 = ~n35684 & n35749;
  assign n35751 = ~n13493 & n32866;
  assign n35752 = ~n14467 & n35751;
  assign n35753 = ~n14573 & n35752;
  assign n35754 = ~n15156 & n35753;
  assign n35755 = n15166 & n35754;
  assign n35756 = ~n13579 & n32871;
  assign n35757 = ~n14467 & n35756;
  assign n35758 = n14574 & n35757;
  assign n35759 = ~n15270 & n35758;
  assign n35760 = n15276 & n35759;
  assign n35761 = n15269 & n35760;
  assign n35762 = ~n35755 & ~n35761;
  assign n35763 = n35750 & n35762;
  assign n35764 = ~n12471 & n30386;
  assign n35765 = ~n14467 & n35764;
  assign n35766 = ~n14466 & n35765;
  assign n35767 = n14574 & n35766;
  assign n35768 = n15599 & n35767;
  assign n35769 = n15595 & n35768;
  assign n35770 = n15593 & n35769;
  assign n35771 = n15615 & n35770;
  assign n35772 = ~n11611 & n32772;
  assign n35773 = ~n14467 & n35772;
  assign n35774 = ~n13820 & n35773;
  assign n35775 = ~n14454 & n35774;
  assign n35776 = ~n14455 & n35775;
  assign n35777 = n14738 & n35776;
  assign n35778 = n14730 & n35777;
  assign n35779 = n14723 & n35778;
  assign n35780 = ~n35771 & ~n35779;
  assign n35781 = n35763 & n35780;
  assign n35782 = n35680 & n35781;
  assign n35783 = n35658 & n35782;
  assign n35784 = n14981 & n22614;
  assign n35785 = ~n3066 & n35784;
  assign n35786 = ~n3983 & n35785;
  assign n35787 = ~n4003 & n35786;
  assign n35788 = ~n4024 & n35787;
  assign n35789 = ~n4999 & n35788;
  assign n35790 = ~n5827 & n35789;
  assign n35791 = ~n6893 & n35790;
  assign n35792 = ~n7890 & n35791;
  assign n35793 = ~n9131 & n35792;
  assign n35794 = ~n14797 & n35793;
  assign n35795 = ~n14796 & n35794;
  assign n35796 = ~n10278 & n35795;
  assign n35797 = ~n11662 & n35796;
  assign n35798 = ~n14795 & n35797;
  assign n35799 = ~n14794 & n35798;
  assign n35800 = n14817 & n35799;
  assign n35801 = n14820 & n35800;
  assign n35802 = n14824 & n35801;
  assign n35803 = n14793 & n35802;
  assign n35804 = n14847 & n35803;
  assign n35805 = n15247 & n32989;
  assign n35806 = ~n5808 & n35805;
  assign n35807 = ~n6056 & n35806;
  assign n35808 = ~n7073 & n35807;
  assign n35809 = ~n8179 & n35808;
  assign n35810 = ~n9344 & n35809;
  assign n35811 = ~n15195 & n35810;
  assign n35812 = ~n15194 & n35811;
  assign n35813 = ~n10594 & n35812;
  assign n35814 = ~n12005 & n35813;
  assign n35815 = ~n14467 & n35814;
  assign n35816 = ~n14572 & n35815;
  assign n35817 = n15208 & n35816;
  assign n35818 = n15211 & n35817;
  assign n35819 = n15215 & n35818;
  assign n35820 = n15193 & n35819;
  assign n35821 = n15238 & n35820;
  assign n35822 = pi188 & ~n9913;
  assign n35823 = n15548 & n35822;
  assign n35824 = ~n9929 & n35823;
  assign n35825 = ~n15497 & n35824;
  assign n35826 = ~n15496 & n35825;
  assign n35827 = ~n11266 & n35826;
  assign n35828 = ~n11588 & n35827;
  assign n35829 = ~n14467 & n35828;
  assign n35830 = ~n14466 & n35829;
  assign n35831 = n14574 & n35830;
  assign n35832 = n15508 & n35831;
  assign n35833 = n15512 & n35832;
  assign n35834 = n15495 & n35833;
  assign n35835 = n15535 & n35834;
  assign n35836 = ~n35821 & ~n35835;
  assign n35837 = ~n35804 & n35836;
  assign n35838 = pi108 & ~n4401;
  assign n35839 = n13494 & n35838;
  assign n35840 = ~n4817 & n35839;
  assign n35841 = ~n4902 & n35840;
  assign n35842 = ~n6001 & n35841;
  assign n35843 = ~n7014 & n35842;
  assign n35844 = ~n8114 & n35843;
  assign n35845 = ~n9276 & n35844;
  assign n35846 = ~n15107 & n35845;
  assign n35847 = ~n15106 & n35846;
  assign n35848 = ~n10523 & n35847;
  assign n35849 = ~n11928 & n35848;
  assign n35850 = ~n14467 & n35849;
  assign n35851 = ~n14573 & n35850;
  assign n35852 = n15122 & n35851;
  assign n35853 = n15125 & n35852;
  assign n35854 = n15129 & n35853;
  assign n35855 = n15105 & n35854;
  assign n35856 = n15152 & n35855;
  assign n35857 = pi236 & ~n14416;
  assign n35858 = n15890 & n35857;
  assign n35859 = ~n14519 & n35858;
  assign n35860 = ~n15742 & n35859;
  assign n35861 = ~n14467 & n35860;
  assign n35862 = ~n14466 & n35861;
  assign n35863 = n14574 & n35862;
  assign n35864 = ~n14577 & n35863;
  assign n35865 = n15756 & n35864;
  assign n35866 = n14457 & n35865;
  assign n35867 = n15854 & n35866;
  assign n35868 = ~n35856 & ~n35867;
  assign n35869 = ~n14467 & n32925;
  assign n35870 = ~n14466 & n35869;
  assign n35871 = n14574 & n35870;
  assign n35872 = n15859 & n35871;
  assign n35873 = n15862 & n35872;
  assign n35874 = n15595 & n35873;
  assign n35875 = n15885 & n35874;
  assign n35876 = n15424 & n24206;
  assign n35877 = ~n7869 & n35876;
  assign n35878 = ~n8346 & n35877;
  assign n35879 = ~n9485 & n35878;
  assign n35880 = ~n15345 & n35879;
  assign n35881 = ~n15344 & n35880;
  assign n35882 = ~n10741 & n35881;
  assign n35883 = ~n12158 & n35882;
  assign n35884 = ~n14467 & n35883;
  assign n35885 = ~n14466 & n35884;
  assign n35886 = n14574 & n35885;
  assign n35887 = n15357 & n35886;
  assign n35888 = n15361 & n35887;
  assign n35889 = n15343 & n35888;
  assign n35890 = n15384 & n35889;
  assign n35891 = ~n35875 & ~n35890;
  assign n35892 = n35868 & n35891;
  assign n35893 = n13408 & n28036;
  assign n35894 = ~n3940 & n35893;
  assign n35895 = ~n4001 & n35894;
  assign n35896 = ~n5043 & n35895;
  assign n35897 = ~n5943 & n35896;
  assign n35898 = ~n6951 & n35897;
  assign n35899 = ~n8037 & n35898;
  assign n35900 = ~n9200 & n35899;
  assign n35901 = ~n15012 & n35900;
  assign n35902 = ~n15011 & n35901;
  assign n35903 = ~n10445 & n35902;
  assign n35904 = ~n11846 & n35903;
  assign n35905 = ~n14467 & n35904;
  assign n35906 = ~n15010 & n35905;
  assign n35907 = n15030 & n35906;
  assign n35908 = n15033 & n35907;
  assign n35909 = n15037 & n35908;
  assign n35910 = n15009 & n35909;
  assign n35911 = n15060 & n35910;
  assign n35912 = n14858 & n27997;
  assign n35913 = ~n1372 & n35912;
  assign n35914 = ~n2243 & n35913;
  assign n35915 = ~n3104 & n35914;
  assign n35916 = ~n3971 & n35915;
  assign n35917 = ~n4003 & n35916;
  assign n35918 = ~n4872 & n35917;
  assign n35919 = ~n5801 & n35918;
  assign n35920 = ~n6739 & n35919;
  assign n35921 = ~n7807 & n35920;
  assign n35922 = ~n8989 & n35921;
  assign n35923 = ~n10273 & n35922;
  assign n35924 = ~n14857 & n35923;
  assign n35925 = ~n14856 & n35924;
  assign n35926 = ~n11499 & n35925;
  assign n35927 = ~n13076 & n35926;
  assign n35928 = ~n14855 & n35927;
  assign n35929 = ~n14854 & n35928;
  assign n35930 = n14879 & n35929;
  assign n35931 = n14882 & n35930;
  assign n35932 = n14886 & n35931;
  assign n35933 = n14853 & n35932;
  assign n35934 = n14909 & n35933;
  assign n35935 = ~n35911 & ~n35934;
  assign n35936 = n15386 & n28055;
  assign n35937 = ~n6784 & n35936;
  assign n35938 = ~n7158 & n35937;
  assign n35939 = ~n8250 & n35938;
  assign n35940 = ~n9414 & n35939;
  assign n35941 = ~n15287 & n35940;
  assign n35942 = ~n15286 & n35941;
  assign n35943 = ~n10667 & n35942;
  assign n35944 = ~n12083 & n35943;
  assign n35945 = ~n14467 & n35944;
  assign n35946 = ~n14466 & n35945;
  assign n35947 = n14574 & n35946;
  assign n35948 = n15302 & n35947;
  assign n35949 = n15306 & n35948;
  assign n35950 = n15285 & n35949;
  assign n35951 = n15329 & n35950;
  assign n35952 = n14749 & n32974;
  assign n35953 = ~n8834 & n35952;
  assign n35954 = ~n10002 & n35953;
  assign n35955 = ~n14747 & n35954;
  assign n35956 = ~n14746 & n35955;
  assign n35957 = ~n11297 & n35956;
  assign n35958 = ~n12240 & n35957;
  assign n35959 = ~n14467 & n35958;
  assign n35960 = ~n14466 & n35959;
  assign n35961 = n14574 & n35960;
  assign n35962 = n14760 & n35961;
  assign n35963 = n14764 & n35962;
  assign n35964 = n14745 & n35963;
  assign n35965 = n14787 & n35964;
  assign n35966 = ~n35951 & ~n35965;
  assign n35967 = n35935 & n35966;
  assign n35968 = n35892 & n35967;
  assign n35969 = n35837 & n35968;
  assign po133 = ~n35783 | ~n35969;
  assign n35971 = pi061 & ~n1740;
  assign n35972 = n13259 & n35971;
  assign n35973 = ~n2242 & n35972;
  assign n35974 = ~n3095 & n35973;
  assign n35975 = ~n3997 & n35974;
  assign n35976 = ~n4003 & n35975;
  assign n35977 = ~n4837 & n35976;
  assign n35978 = ~n5822 & n35977;
  assign n35979 = ~n6820 & n35978;
  assign n35980 = ~n7785 & n35979;
  assign n35981 = ~n9027 & n35980;
  assign n35982 = ~n10245 & n35981;
  assign n35983 = ~n14919 & n35982;
  assign n35984 = ~n14918 & n35983;
  assign n35985 = ~n11536 & n35984;
  assign n35986 = ~n13036 & n35985;
  assign n35987 = ~n14917 & n35986;
  assign n35988 = ~n14916 & n35987;
  assign n35989 = n14940 & n35988;
  assign n35990 = n14943 & n35989;
  assign n35991 = n14947 & n35990;
  assign n35992 = n14915 & n35991;
  assign n35993 = n14970 & n35992;
  assign n35994 = pi245 & ~n14568;
  assign n35995 = ~n14520 & n35994;
  assign n35996 = ~n14467 & n35995;
  assign n35997 = ~n14466 & n35996;
  assign n35998 = n14574 & n35997;
  assign n35999 = ~n14465 & n35998;
  assign n36000 = n14581 & n35999;
  assign n36001 = n14457 & n36000;
  assign n36002 = n14715 & n36001;
  assign n36003 = ~n35993 & ~n36002;
  assign n36004 = pi205 & ~n11168;
  assign n36005 = n15698 & n36004;
  assign n36006 = ~n11188 & n36005;
  assign n36007 = ~n15620 & n36006;
  assign n36008 = ~n15619 & n36007;
  assign n36009 = ~n12380 & n36008;
  assign n36010 = ~n14467 & n36009;
  assign n36011 = ~n14466 & n36010;
  assign n36012 = n14574 & n36011;
  assign n36013 = n15629 & n36012;
  assign n36014 = n15633 & n36013;
  assign n36015 = n15595 & n36014;
  assign n36016 = n15656 & n36015;
  assign n36017 = pi221 & ~n12841;
  assign n36018 = n12775 & n36017;
  assign n36019 = ~n12902 & n36018;
  assign n36020 = ~n15659 & n36019;
  assign n36021 = ~n15658 & n36020;
  assign n36022 = ~n14467 & n36021;
  assign n36023 = ~n14466 & n36022;
  assign n36024 = n14574 & n36023;
  assign n36025 = n15666 & n36024;
  assign n36026 = n15669 & n36025;
  assign n36027 = n15595 & n36026;
  assign n36028 = n15692 & n36027;
  assign n36029 = ~n36016 & ~n36028;
  assign n36030 = n36003 & n36029;
  assign n36031 = ~n11551 & n33104;
  assign n36032 = ~n14467 & n36031;
  assign n36033 = ~n13906 & n36032;
  assign n36034 = ~n14452 & n36033;
  assign n36035 = n14456 & n36034;
  assign n36036 = n15571 & n36035;
  assign n36037 = n15585 & n36036;
  assign n36038 = ~n12181 & n33089;
  assign n36039 = ~n14467 & n36038;
  assign n36040 = ~n13764 & n36039;
  assign n36041 = ~n14455 & n36040;
  assign n36042 = n14737 & n36041;
  assign n36043 = n15463 & n36042;
  assign n36044 = n15452 & n36043;
  assign n36045 = ~n12121 & n33082;
  assign n36046 = ~n14467 & n36045;
  assign n36047 = ~n13726 & n36046;
  assign n36048 = n14737 & n36047;
  assign n36049 = n15417 & n36048;
  assign n36050 = n15407 & n36049;
  assign n36051 = ~n36044 & ~n36050;
  assign n36052 = ~n36037 & n36051;
  assign n36053 = ~n13407 & n33126;
  assign n36054 = ~n14467 & n36053;
  assign n36055 = ~n15067 & n36054;
  assign n36056 = n15074 & n36055;
  assign n36057 = ~n13318 & n33130;
  assign n36058 = ~n14974 & n36057;
  assign n36059 = n14979 & n36058;
  assign n36060 = pi261 & ~n501;
  assign n36061 = n12872 & n36060;
  assign n36062 = n15973 & n36061;
  assign n36063 = n15980 & n36062;
  assign n36064 = n15972 & n36063;
  assign n36065 = n16005 & n36064;
  assign n36066 = ~n1172 & n36065;
  assign n36067 = ~n996 & n36066;
  assign n36068 = ~n2306 & n36067;
  assign n36069 = ~n500 & n36068;
  assign n36070 = n16011 & n36069;
  assign n36071 = n16014 & n36070;
  assign n36072 = n16017 & n36071;
  assign n36073 = n16038 & n36072;
  assign n36074 = n15963 & n36073;
  assign n36075 = n15954 & n36074;
  assign n36076 = ~n7236 & n36075;
  assign n36077 = ~n6137 & n36076;
  assign n36078 = n6193 & n36077;
  assign n36079 = n6134 & n36078;
  assign n36080 = ~n8867 & n36079;
  assign n36081 = ~n7235 & n36080;
  assign n36082 = n7296 & n36081;
  assign n36083 = n7231 & n36082;
  assign n36084 = ~n10027 & n36083;
  assign n36085 = ~n8866 & n36084;
  assign n36086 = n8898 & n36085;
  assign n36087 = n8863 & n36086;
  assign n36088 = pi253 & ~n501;
  assign n36089 = n12872 & n36088;
  assign n36090 = n15973 & n36089;
  assign n36091 = n16069 & n36090;
  assign n36092 = n16063 & n36091;
  assign n36093 = n16088 & n36092;
  assign n36094 = ~n1172 & n36093;
  assign n36095 = ~n996 & n36094;
  assign n36096 = ~n2306 & n36095;
  assign n36097 = ~n500 & n36096;
  assign n36098 = n16094 & n36097;
  assign n36099 = n16016 & n36098;
  assign n36100 = n16054 & n36099;
  assign n36101 = n16113 & n36100;
  assign n36102 = n16184 & n36101;
  assign n36103 = n16048 & n36102;
  assign n36104 = ~n7236 & n36103;
  assign n36105 = ~n6137 & n36104;
  assign n36106 = n6193 & n36105;
  assign n36107 = n6134 & n36106;
  assign n36108 = ~n8867 & n36107;
  assign n36109 = ~n7235 & n36108;
  assign n36110 = n7296 & n36109;
  assign n36111 = n7231 & n36110;
  assign n36112 = ~n10027 & n36111;
  assign n36113 = ~n8866 & n36112;
  assign n36114 = n8898 & n36113;
  assign n36115 = n8863 & n36114;
  assign n36116 = ~n36087 & ~n36115;
  assign n36117 = ~n10788 & ~n36116;
  assign n36118 = ~n10026 & n36117;
  assign n36119 = n10072 & n36118;
  assign n36120 = n10021 & n36119;
  assign n36121 = ~n36059 & ~n36120;
  assign n36122 = ~n36056 & n36121;
  assign n36123 = ~n13493 & n33191;
  assign n36124 = ~n14467 & n36123;
  assign n36125 = ~n14573 & n36124;
  assign n36126 = ~n15156 & n36125;
  assign n36127 = n15166 & n36126;
  assign n36128 = ~n13579 & n33196;
  assign n36129 = ~n14467 & n36128;
  assign n36130 = n14574 & n36129;
  assign n36131 = ~n15270 & n36130;
  assign n36132 = n15276 & n36131;
  assign n36133 = n15269 & n36132;
  assign n36134 = ~n36127 & ~n36133;
  assign n36135 = n36122 & n36134;
  assign n36136 = ~n12471 & n30687;
  assign n36137 = ~n14467 & n36136;
  assign n36138 = ~n14466 & n36137;
  assign n36139 = n14574 & n36138;
  assign n36140 = n15599 & n36139;
  assign n36141 = n15595 & n36140;
  assign n36142 = n15593 & n36141;
  assign n36143 = n15615 & n36142;
  assign n36144 = ~n11611 & n33097;
  assign n36145 = ~n14467 & n36144;
  assign n36146 = ~n13820 & n36145;
  assign n36147 = ~n14454 & n36146;
  assign n36148 = ~n14455 & n36147;
  assign n36149 = n14738 & n36148;
  assign n36150 = n14730 & n36149;
  assign n36151 = n14723 & n36150;
  assign n36152 = ~n36143 & ~n36151;
  assign n36153 = n36135 & n36152;
  assign n36154 = n36052 & n36153;
  assign n36155 = n36030 & n36154;
  assign n36156 = n14981 & n22781;
  assign n36157 = ~n3066 & n36156;
  assign n36158 = ~n3983 & n36157;
  assign n36159 = ~n4003 & n36158;
  assign n36160 = ~n4024 & n36159;
  assign n36161 = ~n4999 & n36160;
  assign n36162 = ~n5827 & n36161;
  assign n36163 = ~n6893 & n36162;
  assign n36164 = ~n7890 & n36163;
  assign n36165 = ~n9131 & n36164;
  assign n36166 = ~n14797 & n36165;
  assign n36167 = ~n14796 & n36166;
  assign n36168 = ~n10278 & n36167;
  assign n36169 = ~n11662 & n36168;
  assign n36170 = ~n14795 & n36169;
  assign n36171 = ~n14794 & n36170;
  assign n36172 = n14817 & n36171;
  assign n36173 = n14820 & n36172;
  assign n36174 = n14824 & n36173;
  assign n36175 = n14793 & n36174;
  assign n36176 = n14847 & n36175;
  assign n36177 = n15247 & n33314;
  assign n36178 = ~n5808 & n36177;
  assign n36179 = ~n6056 & n36178;
  assign n36180 = ~n7073 & n36179;
  assign n36181 = ~n8179 & n36180;
  assign n36182 = ~n9344 & n36181;
  assign n36183 = ~n15195 & n36182;
  assign n36184 = ~n15194 & n36183;
  assign n36185 = ~n10594 & n36184;
  assign n36186 = ~n12005 & n36185;
  assign n36187 = ~n14467 & n36186;
  assign n36188 = ~n14572 & n36187;
  assign n36189 = n15208 & n36188;
  assign n36190 = n15211 & n36189;
  assign n36191 = n15215 & n36190;
  assign n36192 = n15193 & n36191;
  assign n36193 = n15238 & n36192;
  assign n36194 = pi189 & ~n9913;
  assign n36195 = n15548 & n36194;
  assign n36196 = ~n9929 & n36195;
  assign n36197 = ~n15497 & n36196;
  assign n36198 = ~n15496 & n36197;
  assign n36199 = ~n11266 & n36198;
  assign n36200 = ~n11588 & n36199;
  assign n36201 = ~n14467 & n36200;
  assign n36202 = ~n14466 & n36201;
  assign n36203 = n14574 & n36202;
  assign n36204 = n15508 & n36203;
  assign n36205 = n15512 & n36204;
  assign n36206 = n15495 & n36205;
  assign n36207 = n15535 & n36206;
  assign n36208 = ~n36193 & ~n36207;
  assign n36209 = ~n36176 & n36208;
  assign n36210 = pi109 & ~n4401;
  assign n36211 = n13494 & n36210;
  assign n36212 = ~n4817 & n36211;
  assign n36213 = ~n4902 & n36212;
  assign n36214 = ~n6001 & n36213;
  assign n36215 = ~n7014 & n36214;
  assign n36216 = ~n8114 & n36215;
  assign n36217 = ~n9276 & n36216;
  assign n36218 = ~n15107 & n36217;
  assign n36219 = ~n15106 & n36218;
  assign n36220 = ~n10523 & n36219;
  assign n36221 = ~n11928 & n36220;
  assign n36222 = ~n14467 & n36221;
  assign n36223 = ~n14573 & n36222;
  assign n36224 = n15122 & n36223;
  assign n36225 = n15125 & n36224;
  assign n36226 = n15129 & n36225;
  assign n36227 = n15105 & n36226;
  assign n36228 = n15152 & n36227;
  assign n36229 = pi237 & ~n14416;
  assign n36230 = n15890 & n36229;
  assign n36231 = ~n14519 & n36230;
  assign n36232 = ~n15742 & n36231;
  assign n36233 = ~n14467 & n36232;
  assign n36234 = ~n14466 & n36233;
  assign n36235 = n14574 & n36234;
  assign n36236 = ~n14577 & n36235;
  assign n36237 = n15756 & n36236;
  assign n36238 = n14457 & n36237;
  assign n36239 = n15854 & n36238;
  assign n36240 = ~n36228 & ~n36239;
  assign n36241 = ~n14467 & n33250;
  assign n36242 = ~n14466 & n36241;
  assign n36243 = n14574 & n36242;
  assign n36244 = n15859 & n36243;
  assign n36245 = n15862 & n36244;
  assign n36246 = n15595 & n36245;
  assign n36247 = n15885 & n36246;
  assign n36248 = n15424 & n24399;
  assign n36249 = ~n7869 & n36248;
  assign n36250 = ~n8346 & n36249;
  assign n36251 = ~n9485 & n36250;
  assign n36252 = ~n15345 & n36251;
  assign n36253 = ~n15344 & n36252;
  assign n36254 = ~n10741 & n36253;
  assign n36255 = ~n12158 & n36254;
  assign n36256 = ~n14467 & n36255;
  assign n36257 = ~n14466 & n36256;
  assign n36258 = n14574 & n36257;
  assign n36259 = n15357 & n36258;
  assign n36260 = n15361 & n36259;
  assign n36261 = n15343 & n36260;
  assign n36262 = n15384 & n36261;
  assign n36263 = ~n36247 & ~n36262;
  assign n36264 = n36240 & n36263;
  assign n36265 = n13408 & n28302;
  assign n36266 = ~n3940 & n36265;
  assign n36267 = ~n4001 & n36266;
  assign n36268 = ~n5043 & n36267;
  assign n36269 = ~n5943 & n36268;
  assign n36270 = ~n6951 & n36269;
  assign n36271 = ~n8037 & n36270;
  assign n36272 = ~n9200 & n36271;
  assign n36273 = ~n15012 & n36272;
  assign n36274 = ~n15011 & n36273;
  assign n36275 = ~n10445 & n36274;
  assign n36276 = ~n11846 & n36275;
  assign n36277 = ~n14467 & n36276;
  assign n36278 = ~n15010 & n36277;
  assign n36279 = n15030 & n36278;
  assign n36280 = n15033 & n36279;
  assign n36281 = n15037 & n36280;
  assign n36282 = n15009 & n36281;
  assign n36283 = n15060 & n36282;
  assign n36284 = n14858 & n28263;
  assign n36285 = ~n1372 & n36284;
  assign n36286 = ~n2243 & n36285;
  assign n36287 = ~n3104 & n36286;
  assign n36288 = ~n3971 & n36287;
  assign n36289 = ~n4003 & n36288;
  assign n36290 = ~n4872 & n36289;
  assign n36291 = ~n5801 & n36290;
  assign n36292 = ~n6739 & n36291;
  assign n36293 = ~n7807 & n36292;
  assign n36294 = ~n8989 & n36293;
  assign n36295 = ~n10273 & n36294;
  assign n36296 = ~n14857 & n36295;
  assign n36297 = ~n14856 & n36296;
  assign n36298 = ~n11499 & n36297;
  assign n36299 = ~n13076 & n36298;
  assign n36300 = ~n14855 & n36299;
  assign n36301 = ~n14854 & n36300;
  assign n36302 = n14879 & n36301;
  assign n36303 = n14882 & n36302;
  assign n36304 = n14886 & n36303;
  assign n36305 = n14853 & n36304;
  assign n36306 = n14909 & n36305;
  assign n36307 = ~n36283 & ~n36306;
  assign n36308 = n15386 & n28321;
  assign n36309 = ~n6784 & n36308;
  assign n36310 = ~n7158 & n36309;
  assign n36311 = ~n8250 & n36310;
  assign n36312 = ~n9414 & n36311;
  assign n36313 = ~n15287 & n36312;
  assign n36314 = ~n15286 & n36313;
  assign n36315 = ~n10667 & n36314;
  assign n36316 = ~n12083 & n36315;
  assign n36317 = ~n14467 & n36316;
  assign n36318 = ~n14466 & n36317;
  assign n36319 = n14574 & n36318;
  assign n36320 = n15302 & n36319;
  assign n36321 = n15306 & n36320;
  assign n36322 = n15285 & n36321;
  assign n36323 = n15329 & n36322;
  assign n36324 = n14749 & n33299;
  assign n36325 = ~n8834 & n36324;
  assign n36326 = ~n10002 & n36325;
  assign n36327 = ~n14747 & n36326;
  assign n36328 = ~n14746 & n36327;
  assign n36329 = ~n11297 & n36328;
  assign n36330 = ~n12240 & n36329;
  assign n36331 = ~n14467 & n36330;
  assign n36332 = ~n14466 & n36331;
  assign n36333 = n14574 & n36332;
  assign n36334 = n14760 & n36333;
  assign n36335 = n14764 & n36334;
  assign n36336 = n14745 & n36335;
  assign n36337 = n14787 & n36336;
  assign n36338 = ~n36323 & ~n36337;
  assign n36339 = n36307 & n36338;
  assign n36340 = n36264 & n36339;
  assign n36341 = n36209 & n36340;
  assign po134 = ~n36155 | ~n36341;
  assign n36343 = pi062 & ~n1740;
  assign n36344 = n13259 & n36343;
  assign n36345 = ~n2242 & n36344;
  assign n36346 = ~n3095 & n36345;
  assign n36347 = ~n3997 & n36346;
  assign n36348 = ~n4003 & n36347;
  assign n36349 = ~n4837 & n36348;
  assign n36350 = ~n5822 & n36349;
  assign n36351 = ~n6820 & n36350;
  assign n36352 = ~n7785 & n36351;
  assign n36353 = ~n9027 & n36352;
  assign n36354 = ~n10245 & n36353;
  assign n36355 = ~n14919 & n36354;
  assign n36356 = ~n14918 & n36355;
  assign n36357 = ~n11536 & n36356;
  assign n36358 = ~n13036 & n36357;
  assign n36359 = ~n14917 & n36358;
  assign n36360 = ~n14916 & n36359;
  assign n36361 = n14940 & n36360;
  assign n36362 = n14943 & n36361;
  assign n36363 = n14947 & n36362;
  assign n36364 = n14915 & n36363;
  assign n36365 = n14970 & n36364;
  assign n36366 = pi246 & ~n14568;
  assign n36367 = ~n14520 & n36366;
  assign n36368 = ~n14467 & n36367;
  assign n36369 = ~n14466 & n36368;
  assign n36370 = n14574 & n36369;
  assign n36371 = ~n14465 & n36370;
  assign n36372 = n14581 & n36371;
  assign n36373 = n14457 & n36372;
  assign n36374 = n14715 & n36373;
  assign n36375 = ~n36365 & ~n36374;
  assign n36376 = pi206 & ~n11168;
  assign n36377 = n15698 & n36376;
  assign n36378 = ~n11188 & n36377;
  assign n36379 = ~n15620 & n36378;
  assign n36380 = ~n15619 & n36379;
  assign n36381 = ~n12380 & n36380;
  assign n36382 = ~n14467 & n36381;
  assign n36383 = ~n14466 & n36382;
  assign n36384 = n14574 & n36383;
  assign n36385 = n15629 & n36384;
  assign n36386 = n15633 & n36385;
  assign n36387 = n15595 & n36386;
  assign n36388 = n15656 & n36387;
  assign n36389 = pi222 & ~n12841;
  assign n36390 = n12775 & n36389;
  assign n36391 = ~n12902 & n36390;
  assign n36392 = ~n15659 & n36391;
  assign n36393 = ~n15658 & n36392;
  assign n36394 = ~n14467 & n36393;
  assign n36395 = ~n14466 & n36394;
  assign n36396 = n14574 & n36395;
  assign n36397 = n15666 & n36396;
  assign n36398 = n15669 & n36397;
  assign n36399 = n15595 & n36398;
  assign n36400 = n15692 & n36399;
  assign n36401 = ~n36388 & ~n36400;
  assign n36402 = n36375 & n36401;
  assign n36403 = ~n11551 & n33429;
  assign n36404 = ~n14467 & n36403;
  assign n36405 = ~n13906 & n36404;
  assign n36406 = ~n14452 & n36405;
  assign n36407 = n14456 & n36406;
  assign n36408 = n15571 & n36407;
  assign n36409 = n15585 & n36408;
  assign n36410 = ~n12181 & n33414;
  assign n36411 = ~n14467 & n36410;
  assign n36412 = ~n13764 & n36411;
  assign n36413 = ~n14455 & n36412;
  assign n36414 = n14737 & n36413;
  assign n36415 = n15463 & n36414;
  assign n36416 = n15452 & n36415;
  assign n36417 = ~n12121 & n33407;
  assign n36418 = ~n14467 & n36417;
  assign n36419 = ~n13726 & n36418;
  assign n36420 = n14737 & n36419;
  assign n36421 = n15417 & n36420;
  assign n36422 = n15407 & n36421;
  assign n36423 = ~n36416 & ~n36422;
  assign n36424 = ~n36409 & n36423;
  assign n36425 = ~n13407 & n33451;
  assign n36426 = ~n14467 & n36425;
  assign n36427 = ~n15067 & n36426;
  assign n36428 = n15074 & n36427;
  assign n36429 = ~n13318 & n33455;
  assign n36430 = ~n14974 & n36429;
  assign n36431 = n14979 & n36430;
  assign n36432 = pi262 & ~n501;
  assign n36433 = n12872 & n36432;
  assign n36434 = n15973 & n36433;
  assign n36435 = n15980 & n36434;
  assign n36436 = n15972 & n36435;
  assign n36437 = n16005 & n36436;
  assign n36438 = ~n1172 & n36437;
  assign n36439 = ~n996 & n36438;
  assign n36440 = ~n2306 & n36439;
  assign n36441 = ~n500 & n36440;
  assign n36442 = n16011 & n36441;
  assign n36443 = n16014 & n36442;
  assign n36444 = n16017 & n36443;
  assign n36445 = n16038 & n36444;
  assign n36446 = n15963 & n36445;
  assign n36447 = n15954 & n36446;
  assign n36448 = ~n7236 & n36447;
  assign n36449 = ~n6137 & n36448;
  assign n36450 = n6193 & n36449;
  assign n36451 = n6134 & n36450;
  assign n36452 = ~n8867 & n36451;
  assign n36453 = ~n7235 & n36452;
  assign n36454 = n7296 & n36453;
  assign n36455 = n7231 & n36454;
  assign n36456 = ~n10027 & n36455;
  assign n36457 = ~n8866 & n36456;
  assign n36458 = n8898 & n36457;
  assign n36459 = n8863 & n36458;
  assign n36460 = pi254 & ~n501;
  assign n36461 = n12872 & n36460;
  assign n36462 = n15973 & n36461;
  assign n36463 = n16069 & n36462;
  assign n36464 = n16063 & n36463;
  assign n36465 = n16088 & n36464;
  assign n36466 = ~n1172 & n36465;
  assign n36467 = ~n996 & n36466;
  assign n36468 = ~n2306 & n36467;
  assign n36469 = ~n500 & n36468;
  assign n36470 = n16094 & n36469;
  assign n36471 = n16016 & n36470;
  assign n36472 = n16054 & n36471;
  assign n36473 = n16113 & n36472;
  assign n36474 = n16184 & n36473;
  assign n36475 = n16048 & n36474;
  assign n36476 = ~n7236 & n36475;
  assign n36477 = ~n6137 & n36476;
  assign n36478 = n6193 & n36477;
  assign n36479 = n6134 & n36478;
  assign n36480 = ~n8867 & n36479;
  assign n36481 = ~n7235 & n36480;
  assign n36482 = n7296 & n36481;
  assign n36483 = n7231 & n36482;
  assign n36484 = ~n10027 & n36483;
  assign n36485 = ~n8866 & n36484;
  assign n36486 = n8898 & n36485;
  assign n36487 = n8863 & n36486;
  assign n36488 = ~n36459 & ~n36487;
  assign n36489 = ~n10788 & ~n36488;
  assign n36490 = ~n10026 & n36489;
  assign n36491 = n10072 & n36490;
  assign n36492 = n10021 & n36491;
  assign n36493 = ~n36431 & ~n36492;
  assign n36494 = ~n36428 & n36493;
  assign n36495 = ~n13493 & n33516;
  assign n36496 = ~n14467 & n36495;
  assign n36497 = ~n14573 & n36496;
  assign n36498 = ~n15156 & n36497;
  assign n36499 = n15166 & n36498;
  assign n36500 = ~n13579 & n33521;
  assign n36501 = ~n14467 & n36500;
  assign n36502 = n14574 & n36501;
  assign n36503 = ~n15270 & n36502;
  assign n36504 = n15276 & n36503;
  assign n36505 = n15269 & n36504;
  assign n36506 = ~n36499 & ~n36505;
  assign n36507 = n36494 & n36506;
  assign n36508 = ~n12471 & n30988;
  assign n36509 = ~n14467 & n36508;
  assign n36510 = ~n14466 & n36509;
  assign n36511 = n14574 & n36510;
  assign n36512 = n15599 & n36511;
  assign n36513 = n15595 & n36512;
  assign n36514 = n15593 & n36513;
  assign n36515 = n15615 & n36514;
  assign n36516 = ~n11611 & n33422;
  assign n36517 = ~n14467 & n36516;
  assign n36518 = ~n13820 & n36517;
  assign n36519 = ~n14454 & n36518;
  assign n36520 = ~n14455 & n36519;
  assign n36521 = n14738 & n36520;
  assign n36522 = n14730 & n36521;
  assign n36523 = n14723 & n36522;
  assign n36524 = ~n36515 & ~n36523;
  assign n36525 = n36507 & n36524;
  assign n36526 = n36424 & n36525;
  assign n36527 = n36402 & n36526;
  assign n36528 = n14981 & n22948;
  assign n36529 = ~n3066 & n36528;
  assign n36530 = ~n3983 & n36529;
  assign n36531 = ~n4003 & n36530;
  assign n36532 = ~n4024 & n36531;
  assign n36533 = ~n4999 & n36532;
  assign n36534 = ~n5827 & n36533;
  assign n36535 = ~n6893 & n36534;
  assign n36536 = ~n7890 & n36535;
  assign n36537 = ~n9131 & n36536;
  assign n36538 = ~n14797 & n36537;
  assign n36539 = ~n14796 & n36538;
  assign n36540 = ~n10278 & n36539;
  assign n36541 = ~n11662 & n36540;
  assign n36542 = ~n14795 & n36541;
  assign n36543 = ~n14794 & n36542;
  assign n36544 = n14817 & n36543;
  assign n36545 = n14820 & n36544;
  assign n36546 = n14824 & n36545;
  assign n36547 = n14793 & n36546;
  assign n36548 = n14847 & n36547;
  assign n36549 = n15247 & n33639;
  assign n36550 = ~n5808 & n36549;
  assign n36551 = ~n6056 & n36550;
  assign n36552 = ~n7073 & n36551;
  assign n36553 = ~n8179 & n36552;
  assign n36554 = ~n9344 & n36553;
  assign n36555 = ~n15195 & n36554;
  assign n36556 = ~n15194 & n36555;
  assign n36557 = ~n10594 & n36556;
  assign n36558 = ~n12005 & n36557;
  assign n36559 = ~n14467 & n36558;
  assign n36560 = ~n14572 & n36559;
  assign n36561 = n15208 & n36560;
  assign n36562 = n15211 & n36561;
  assign n36563 = n15215 & n36562;
  assign n36564 = n15193 & n36563;
  assign n36565 = n15238 & n36564;
  assign n36566 = pi190 & ~n9913;
  assign n36567 = n15548 & n36566;
  assign n36568 = ~n9929 & n36567;
  assign n36569 = ~n15497 & n36568;
  assign n36570 = ~n15496 & n36569;
  assign n36571 = ~n11266 & n36570;
  assign n36572 = ~n11588 & n36571;
  assign n36573 = ~n14467 & n36572;
  assign n36574 = ~n14466 & n36573;
  assign n36575 = n14574 & n36574;
  assign n36576 = n15508 & n36575;
  assign n36577 = n15512 & n36576;
  assign n36578 = n15495 & n36577;
  assign n36579 = n15535 & n36578;
  assign n36580 = ~n36565 & ~n36579;
  assign n36581 = ~n36548 & n36580;
  assign n36582 = pi110 & ~n4401;
  assign n36583 = n13494 & n36582;
  assign n36584 = ~n4817 & n36583;
  assign n36585 = ~n4902 & n36584;
  assign n36586 = ~n6001 & n36585;
  assign n36587 = ~n7014 & n36586;
  assign n36588 = ~n8114 & n36587;
  assign n36589 = ~n9276 & n36588;
  assign n36590 = ~n15107 & n36589;
  assign n36591 = ~n15106 & n36590;
  assign n36592 = ~n10523 & n36591;
  assign n36593 = ~n11928 & n36592;
  assign n36594 = ~n14467 & n36593;
  assign n36595 = ~n14573 & n36594;
  assign n36596 = n15122 & n36595;
  assign n36597 = n15125 & n36596;
  assign n36598 = n15129 & n36597;
  assign n36599 = n15105 & n36598;
  assign n36600 = n15152 & n36599;
  assign n36601 = pi238 & ~n14416;
  assign n36602 = n15890 & n36601;
  assign n36603 = ~n14519 & n36602;
  assign n36604 = ~n15742 & n36603;
  assign n36605 = ~n14467 & n36604;
  assign n36606 = ~n14466 & n36605;
  assign n36607 = n14574 & n36606;
  assign n36608 = ~n14577 & n36607;
  assign n36609 = n15756 & n36608;
  assign n36610 = n14457 & n36609;
  assign n36611 = n15854 & n36610;
  assign n36612 = ~n36600 & ~n36611;
  assign n36613 = ~n14467 & n33575;
  assign n36614 = ~n14466 & n36613;
  assign n36615 = n14574 & n36614;
  assign n36616 = n15859 & n36615;
  assign n36617 = n15862 & n36616;
  assign n36618 = n15595 & n36617;
  assign n36619 = n15885 & n36618;
  assign n36620 = n15424 & n24592;
  assign n36621 = ~n7869 & n36620;
  assign n36622 = ~n8346 & n36621;
  assign n36623 = ~n9485 & n36622;
  assign n36624 = ~n15345 & n36623;
  assign n36625 = ~n15344 & n36624;
  assign n36626 = ~n10741 & n36625;
  assign n36627 = ~n12158 & n36626;
  assign n36628 = ~n14467 & n36627;
  assign n36629 = ~n14466 & n36628;
  assign n36630 = n14574 & n36629;
  assign n36631 = n15357 & n36630;
  assign n36632 = n15361 & n36631;
  assign n36633 = n15343 & n36632;
  assign n36634 = n15384 & n36633;
  assign n36635 = ~n36619 & ~n36634;
  assign n36636 = n36612 & n36635;
  assign n36637 = n13408 & n28568;
  assign n36638 = ~n3940 & n36637;
  assign n36639 = ~n4001 & n36638;
  assign n36640 = ~n5043 & n36639;
  assign n36641 = ~n5943 & n36640;
  assign n36642 = ~n6951 & n36641;
  assign n36643 = ~n8037 & n36642;
  assign n36644 = ~n9200 & n36643;
  assign n36645 = ~n15012 & n36644;
  assign n36646 = ~n15011 & n36645;
  assign n36647 = ~n10445 & n36646;
  assign n36648 = ~n11846 & n36647;
  assign n36649 = ~n14467 & n36648;
  assign n36650 = ~n15010 & n36649;
  assign n36651 = n15030 & n36650;
  assign n36652 = n15033 & n36651;
  assign n36653 = n15037 & n36652;
  assign n36654 = n15009 & n36653;
  assign n36655 = n15060 & n36654;
  assign n36656 = n14858 & n28529;
  assign n36657 = ~n1372 & n36656;
  assign n36658 = ~n2243 & n36657;
  assign n36659 = ~n3104 & n36658;
  assign n36660 = ~n3971 & n36659;
  assign n36661 = ~n4003 & n36660;
  assign n36662 = ~n4872 & n36661;
  assign n36663 = ~n5801 & n36662;
  assign n36664 = ~n6739 & n36663;
  assign n36665 = ~n7807 & n36664;
  assign n36666 = ~n8989 & n36665;
  assign n36667 = ~n10273 & n36666;
  assign n36668 = ~n14857 & n36667;
  assign n36669 = ~n14856 & n36668;
  assign n36670 = ~n11499 & n36669;
  assign n36671 = ~n13076 & n36670;
  assign n36672 = ~n14855 & n36671;
  assign n36673 = ~n14854 & n36672;
  assign n36674 = n14879 & n36673;
  assign n36675 = n14882 & n36674;
  assign n36676 = n14886 & n36675;
  assign n36677 = n14853 & n36676;
  assign n36678 = n14909 & n36677;
  assign n36679 = ~n36655 & ~n36678;
  assign n36680 = n15386 & n28587;
  assign n36681 = ~n6784 & n36680;
  assign n36682 = ~n7158 & n36681;
  assign n36683 = ~n8250 & n36682;
  assign n36684 = ~n9414 & n36683;
  assign n36685 = ~n15287 & n36684;
  assign n36686 = ~n15286 & n36685;
  assign n36687 = ~n10667 & n36686;
  assign n36688 = ~n12083 & n36687;
  assign n36689 = ~n14467 & n36688;
  assign n36690 = ~n14466 & n36689;
  assign n36691 = n14574 & n36690;
  assign n36692 = n15302 & n36691;
  assign n36693 = n15306 & n36692;
  assign n36694 = n15285 & n36693;
  assign n36695 = n15329 & n36694;
  assign n36696 = n14749 & n33624;
  assign n36697 = ~n8834 & n36696;
  assign n36698 = ~n10002 & n36697;
  assign n36699 = ~n14747 & n36698;
  assign n36700 = ~n14746 & n36699;
  assign n36701 = ~n11297 & n36700;
  assign n36702 = ~n12240 & n36701;
  assign n36703 = ~n14467 & n36702;
  assign n36704 = ~n14466 & n36703;
  assign n36705 = n14574 & n36704;
  assign n36706 = n14760 & n36705;
  assign n36707 = n14764 & n36706;
  assign n36708 = n14745 & n36707;
  assign n36709 = n14787 & n36708;
  assign n36710 = ~n36695 & ~n36709;
  assign n36711 = n36679 & n36710;
  assign n36712 = n36636 & n36711;
  assign n36713 = n36581 & n36712;
  assign po135 = ~n36527 | ~n36713;
  assign n36715 = pi247 & ~n16144;
  assign n36716 = ~n16175 & n36715;
  assign n36717 = ~n16360 & n36716;
  assign n36718 = ~n17630 & n36717;
  assign n36719 = ~n16216 & n36718;
  assign n36720 = ~n16215 & n36719;
  assign n36721 = n16222 & n36720;
  assign n36722 = n17637 & n36721;
  assign n36723 = n17629 & n36722;
  assign n36724 = n17628 & n36723;
  assign n36725 = n17736 & n36724;
  assign n36726 = pi087 & ~n3710;
  assign n36727 = ~n3650 & n36726;
  assign n36728 = ~n3940 & n36727;
  assign n36729 = ~n4001 & n36728;
  assign n36730 = ~n5043 & n36729;
  assign n36731 = ~n5943 & n36730;
  assign n36732 = ~n6951 & n36731;
  assign n36733 = ~n8037 & n36732;
  assign n36734 = ~n9200 & n36733;
  assign n36735 = ~n16555 & n36734;
  assign n36736 = ~n16554 & n36735;
  assign n36737 = ~n10445 & n36736;
  assign n36738 = ~n11846 & n36737;
  assign n36739 = ~n13393 & n36738;
  assign n36740 = ~n16216 & n36739;
  assign n36741 = ~n16553 & n36740;
  assign n36742 = n16573 & n36741;
  assign n36743 = n16576 & n36742;
  assign n36744 = n16580 & n36743;
  assign n36745 = n16552 & n36744;
  assign n36746 = n16605 & n36745;
  assign n36747 = ~n36725 & ~n36746;
  assign n36748 = pi183 & ~n9913;
  assign n36749 = ~n9763 & n36748;
  assign n36750 = ~n9929 & n36749;
  assign n36751 = ~n17263 & n36750;
  assign n36752 = ~n17262 & n36751;
  assign n36753 = ~n11266 & n36752;
  assign n36754 = ~n11588 & n36753;
  assign n36755 = ~n13859 & n36754;
  assign n36756 = ~n16216 & n36755;
  assign n36757 = ~n16215 & n36756;
  assign n36758 = n16222 & n36757;
  assign n36759 = n17273 & n36758;
  assign n36760 = n17277 & n36759;
  assign n36761 = n17261 & n36760;
  assign n36762 = n17302 & n36761;
  assign n36763 = pi215 & ~n12743;
  assign n36764 = ~n12773 & n36763;
  assign n36765 = ~n12902 & n36764;
  assign n36766 = ~n17419 & n36765;
  assign n36767 = ~n17418 & n36766;
  assign n36768 = ~n14009 & n36767;
  assign n36769 = ~n16216 & n36768;
  assign n36770 = ~n16215 & n36769;
  assign n36771 = n16222 & n36770;
  assign n36772 = n17427 & n36771;
  assign n36773 = n17431 & n36772;
  assign n36774 = n16214 & n36773;
  assign n36775 = n17456 & n36774;
  assign n36776 = ~n36762 & ~n36775;
  assign n36777 = n36747 & n36776;
  assign n36778 = ~n13764 & n33907;
  assign n36779 = ~n16216 & n36778;
  assign n36780 = ~n15465 & n36779;
  assign n36781 = ~n16209 & n36780;
  assign n36782 = n17086 & n36781;
  assign n36783 = n17133 & n36782;
  assign n36784 = n17122 & n36783;
  assign n36785 = ~n13726 & n33808;
  assign n36786 = ~n16216 & n36785;
  assign n36787 = ~n15419 & n36786;
  assign n36788 = n17086 & n36787;
  assign n36789 = n17094 & n36788;
  assign n36790 = n17083 & n36789;
  assign n36791 = ~n36784 & ~n36790;
  assign n36792 = ~n13093 & n31309;
  assign n36793 = ~n16216 & n36792;
  assign n36794 = ~n16215 & n36793;
  assign n36795 = n16222 & n36794;
  assign n36796 = n17516 & n36795;
  assign n36797 = n16214 & n36796;
  assign n36798 = n17512 & n36797;
  assign n36799 = n17534 & n36798;
  assign n36800 = ~n14073 & n33800;
  assign n36801 = ~n16216 & n36800;
  assign n36802 = ~n15616 & n36801;
  assign n36803 = ~n16224 & n36802;
  assign n36804 = n17086 & n36803;
  assign n36805 = n17351 & n36804;
  assign n36806 = n17350 & n36805;
  assign n36807 = n17370 & n36806;
  assign n36808 = ~n36799 & ~n36807;
  assign n36809 = n36791 & n36808;
  assign n36810 = ~n15075 & n33824;
  assign n36811 = ~n16216 & n36810;
  assign n36812 = ~n16537 & n36811;
  assign n36813 = n16544 & n36812;
  assign n36814 = ~n16831 & n33828;
  assign n36815 = ~n16829 & n36814;
  assign n36816 = n16836 & n36815;
  assign n36817 = pi263 & ~n501;
  assign n36818 = n12872 & n36817;
  assign n36819 = n17949 & n36818;
  assign n36820 = n17954 & n36819;
  assign n36821 = n17947 & n36820;
  assign n36822 = n17982 & n36821;
  assign n36823 = ~n1172 & n36822;
  assign n36824 = ~n996 & n36823;
  assign n36825 = ~n2306 & n36824;
  assign n36826 = ~n500 & n36825;
  assign n36827 = n17940 & n36826;
  assign n36828 = n17991 & n36827;
  assign n36829 = n17938 & n36828;
  assign n36830 = n17929 & n36829;
  assign n36831 = n17921 & n36830;
  assign n36832 = n18029 & n36831;
  assign n36833 = ~n7236 & n36832;
  assign n36834 = ~n6137 & n36833;
  assign n36835 = n6193 & n36834;
  assign n36836 = n6134 & n36835;
  assign n36837 = ~n8867 & n36836;
  assign n36838 = ~n7235 & n36837;
  assign n36839 = n7296 & n36838;
  assign n36840 = n7231 & n36839;
  assign n36841 = ~n10027 & n36840;
  assign n36842 = ~n8866 & n36841;
  assign n36843 = n8898 & n36842;
  assign n36844 = n8863 & n36843;
  assign n36845 = pi271 & ~n501;
  assign n36846 = n12872 & n36845;
  assign n36847 = n18049 & n36846;
  assign n36848 = n18053 & n36847;
  assign n36849 = n18047 & n36848;
  assign n36850 = n18080 & n36849;
  assign n36851 = ~n1172 & n36850;
  assign n36852 = ~n996 & n36851;
  assign n36853 = ~n2306 & n36852;
  assign n36854 = ~n500 & n36853;
  assign n36855 = n18038 & n36854;
  assign n36856 = n18037 & n36855;
  assign n36857 = n18088 & n36856;
  assign n36858 = n18106 & n36857;
  assign n36859 = n18035 & n36858;
  assign n36860 = n18134 & n36859;
  assign n36861 = ~n7236 & n36860;
  assign n36862 = ~n6137 & n36861;
  assign n36863 = n6193 & n36862;
  assign n36864 = n6134 & n36863;
  assign n36865 = ~n8867 & n36864;
  assign n36866 = ~n7235 & n36865;
  assign n36867 = n7296 & n36866;
  assign n36868 = n7231 & n36867;
  assign n36869 = ~n10027 & n36868;
  assign n36870 = ~n8866 & n36869;
  assign n36871 = n8898 & n36870;
  assign n36872 = n8863 & n36871;
  assign n36873 = ~n36844 & ~n36872;
  assign n36874 = ~n10788 & ~n36873;
  assign n36875 = ~n10026 & n36874;
  assign n36876 = n10072 & n36875;
  assign n36877 = n10021 & n36876;
  assign n36878 = ~n36816 & ~n36877;
  assign n36879 = ~n36813 & n36878;
  assign n36880 = ~n15278 & n33894;
  assign n36881 = ~n16216 & n36880;
  assign n36882 = n16939 & n36881;
  assign n36883 = ~n16937 & n36882;
  assign n36884 = n16944 & n36883;
  assign n36885 = n16936 & n36884;
  assign n36886 = ~n15167 & n33900;
  assign n36887 = ~n16216 & n36886;
  assign n36888 = ~n16220 & n36887;
  assign n36889 = ~n16466 & n36888;
  assign n36890 = n16476 & n36889;
  assign n36891 = ~n36885 & ~n36890;
  assign n36892 = n36879 & n36891;
  assign n36893 = ~n13820 & n33814;
  assign n36894 = ~n16216 & n36893;
  assign n36895 = ~n14741 & n36894;
  assign n36896 = ~n16209 & n36895;
  assign n36897 = ~n16211 & n36896;
  assign n36898 = n17238 & n36897;
  assign n36899 = n17232 & n36898;
  assign n36900 = n17225 & n36899;
  assign n36901 = ~n13906 & n33914;
  assign n36902 = ~n16216 & n36901;
  assign n36903 = ~n15586 & n36902;
  assign n36904 = ~n16208 & n36903;
  assign n36905 = n17257 & n36904;
  assign n36906 = n17328 & n36905;
  assign n36907 = n17342 & n36906;
  assign n36908 = ~n36900 & ~n36907;
  assign n36909 = n36892 & n36908;
  assign n36910 = n36809 & n36909;
  assign n36911 = n36777 & n36910;
  assign n36912 = pi119 & ~n5686;
  assign n36913 = ~n5349 & n36912;
  assign n36914 = ~n5808 & n36913;
  assign n36915 = ~n6056 & n36914;
  assign n36916 = ~n7073 & n36915;
  assign n36917 = ~n8179 & n36916;
  assign n36918 = ~n9344 & n36917;
  assign n36919 = ~n16418 & n36918;
  assign n36920 = ~n16361 & n36919;
  assign n36921 = ~n10594 & n36920;
  assign n36922 = ~n12005 & n36921;
  assign n36923 = ~n13558 & n36922;
  assign n36924 = ~n16216 & n36923;
  assign n36925 = ~n16215 & n36924;
  assign n36926 = n16432 & n36925;
  assign n36927 = n16435 & n36926;
  assign n36928 = n16439 & n36927;
  assign n36929 = n16305 & n36928;
  assign n36930 = n16464 & n36929;
  assign n36931 = pi071 & ~n2602;
  assign n36932 = ~n2783 & n36931;
  assign n36933 = ~n3066 & n36932;
  assign n36934 = ~n3983 & n36933;
  assign n36935 = ~n4003 & n36934;
  assign n36936 = ~n4024 & n36935;
  assign n36937 = ~n4999 & n36936;
  assign n36938 = ~n5827 & n36937;
  assign n36939 = ~n6893 & n36938;
  assign n36940 = ~n7890 & n36939;
  assign n36941 = ~n9131 & n36940;
  assign n36942 = ~n16617 & n36941;
  assign n36943 = ~n16616 & n36942;
  assign n36944 = ~n10278 & n36943;
  assign n36945 = ~n11662 & n36944;
  assign n36946 = ~n13191 & n36945;
  assign n36947 = ~n16615 & n36946;
  assign n36948 = ~n16614 & n36947;
  assign n36949 = n16636 & n36948;
  assign n36950 = n16639 & n36949;
  assign n36951 = n16643 & n36950;
  assign n36952 = n16613 & n36951;
  assign n36953 = n16668 & n36952;
  assign n36954 = ~n36930 & ~n36953;
  assign n36955 = pi167 & ~n8633;
  assign n36956 = ~n8455 & n36955;
  assign n36957 = ~n8834 & n36956;
  assign n36958 = ~n10002 & n36957;
  assign n36959 = ~n17152 & n36958;
  assign n36960 = ~n17151 & n36959;
  assign n36961 = ~n11297 & n36960;
  assign n36962 = ~n12240 & n36961;
  assign n36963 = ~n13135 & n36962;
  assign n36964 = ~n16216 & n36963;
  assign n36965 = ~n16215 & n36964;
  assign n36966 = n16222 & n36965;
  assign n36967 = n17163 & n36966;
  assign n36968 = n17167 & n36967;
  assign n36969 = n17150 & n36968;
  assign n36970 = n17192 & n36969;
  assign n36971 = ~n6401 & n31316;
  assign n36972 = ~n6784 & n36971;
  assign n36973 = ~n7158 & n36972;
  assign n36974 = ~n8250 & n36973;
  assign n36975 = ~n9414 & n36974;
  assign n36976 = ~n16957 & n36975;
  assign n36977 = ~n16956 & n36976;
  assign n36978 = ~n10667 & n36977;
  assign n36979 = ~n12083 & n36978;
  assign n36980 = ~n13644 & n36979;
  assign n36981 = ~n16216 & n36980;
  assign n36982 = ~n16215 & n36981;
  assign n36983 = n16222 & n36982;
  assign n36984 = n16971 & n36983;
  assign n36985 = n16975 & n36984;
  assign n36986 = n16955 & n36985;
  assign n36987 = n17000 & n36986;
  assign n36988 = ~n36970 & ~n36987;
  assign n36989 = n36954 & n36988;
  assign n36990 = ~n1372 & n31117;
  assign n36991 = ~n2243 & n36990;
  assign n36992 = ~n3104 & n36991;
  assign n36993 = ~n3971 & n36992;
  assign n36994 = ~n16682 & n36993;
  assign n36995 = ~n4872 & n36994;
  assign n36996 = ~n5801 & n36995;
  assign n36997 = ~n6739 & n36996;
  assign n36998 = ~n7807 & n36997;
  assign n36999 = ~n8989 & n36998;
  assign n37000 = ~n10273 & n36999;
  assign n37001 = ~n16680 & n37000;
  assign n37002 = ~n16679 & n37001;
  assign n37003 = ~n11499 & n37002;
  assign n37004 = ~n13076 & n37003;
  assign n37005 = ~n14698 & n37004;
  assign n37006 = ~n16678 & n37005;
  assign n37007 = ~n16677 & n37006;
  assign n37008 = n16704 & n37007;
  assign n37009 = n16707 & n37008;
  assign n37010 = n16711 & n37009;
  assign n37011 = n16676 & n37010;
  assign n37012 = n16736 & n37011;
  assign n37013 = ~n11042 & n34063;
  assign n37014 = ~n11188 & n37013;
  assign n37015 = ~n17378 & n37014;
  assign n37016 = ~n17377 & n37015;
  assign n37017 = ~n12380 & n37016;
  assign n37018 = ~n14045 & n37017;
  assign n37019 = ~n16216 & n37018;
  assign n37020 = ~n16215 & n37019;
  assign n37021 = n16222 & n37020;
  assign n37022 = n17387 & n37021;
  assign n37023 = n17391 & n37022;
  assign n37024 = n17376 & n37023;
  assign n37025 = n17416 & n37024;
  assign n37026 = ~n37012 & ~n37025;
  assign n37027 = pi103 & ~n4401;
  assign n37028 = ~n4460 & n37027;
  assign n37029 = ~n4817 & n37028;
  assign n37030 = ~n4902 & n37029;
  assign n37031 = ~n6001 & n37030;
  assign n37032 = ~n7014 & n37031;
  assign n37033 = ~n8114 & n37032;
  assign n37034 = ~n9276 & n37033;
  assign n37035 = ~n16486 & n37034;
  assign n37036 = ~n16485 & n37035;
  assign n37037 = ~n10523 & n37036;
  assign n37038 = ~n11928 & n37037;
  assign n37039 = ~n13479 & n37038;
  assign n37040 = ~n16216 & n37039;
  assign n37041 = ~n16220 & n37040;
  assign n37042 = n16503 & n37041;
  assign n37043 = n16506 & n37042;
  assign n37044 = n16510 & n37043;
  assign n37045 = n16484 & n37044;
  assign n37046 = n16535 & n37045;
  assign n37047 = pi055 & ~n1526;
  assign n37048 = ~n1556 & n37047;
  assign n37049 = ~n2242 & n37048;
  assign n37050 = ~n3095 & n37049;
  assign n37051 = ~n3997 & n37050;
  assign n37052 = ~n4003 & n37051;
  assign n37053 = ~n4837 & n37052;
  assign n37054 = ~n5822 & n37053;
  assign n37055 = ~n6820 & n37054;
  assign n37056 = ~n7785 & n37055;
  assign n37057 = ~n9027 & n37056;
  assign n37058 = ~n10245 & n37057;
  assign n37059 = ~n16748 & n37058;
  assign n37060 = ~n16747 & n37059;
  assign n37061 = ~n11536 & n37060;
  assign n37062 = ~n13036 & n37061;
  assign n37063 = ~n14653 & n37062;
  assign n37064 = ~n16746 & n37063;
  assign n37065 = ~n16745 & n37064;
  assign n37066 = n16770 & n37065;
  assign n37067 = n16773 & n37066;
  assign n37068 = n16777 & n37067;
  assign n37069 = n16744 & n37068;
  assign n37070 = n16802 & n37069;
  assign n37071 = ~n37046 & ~n37070;
  assign n37072 = n37026 & n37071;
  assign n37073 = ~n7505 & n34024;
  assign n37074 = ~n7869 & n37073;
  assign n37075 = ~n8346 & n37074;
  assign n37076 = ~n9485 & n37075;
  assign n37077 = ~n17018 & n37076;
  assign n37078 = ~n17017 & n37077;
  assign n37079 = ~n10741 & n37078;
  assign n37080 = ~n12158 & n37079;
  assign n37081 = ~n13693 & n37080;
  assign n37082 = ~n16216 & n37081;
  assign n37083 = ~n16215 & n37082;
  assign n37084 = n16222 & n37083;
  assign n37085 = n17031 & n37084;
  assign n37086 = n17035 & n37085;
  assign n37087 = n17016 & n37086;
  assign n37088 = n17060 & n37087;
  assign n37089 = ~n16216 & n33944;
  assign n37090 = ~n16215 & n37089;
  assign n37091 = n16222 & n37090;
  assign n37092 = n16225 & n37091;
  assign n37093 = n16229 & n37092;
  assign n37094 = n16214 & n37093;
  assign n37095 = n16297 & n37094;
  assign n37096 = ~n37088 & ~n37095;
  assign n37097 = pi231 & ~n14350;
  assign n37098 = ~n14381 & n37097;
  assign n37099 = ~n14519 & n37098;
  assign n37100 = ~n17537 & n37099;
  assign n37101 = ~n17536 & n37100;
  assign n37102 = ~n16216 & n37101;
  assign n37103 = ~n16215 & n37102;
  assign n37104 = n16222 & n37103;
  assign n37105 = n17544 & n37104;
  assign n37106 = n17547 & n37105;
  assign n37107 = n16214 & n37106;
  assign n37108 = n17572 & n37107;
  assign n37109 = pi255 & ~n16417;
  assign n37110 = ~n17766 & n37109;
  assign n37111 = ~n16216 & n37110;
  assign n37112 = ~n16215 & n37111;
  assign n37113 = n16222 & n37112;
  assign n37114 = n17637 & n37113;
  assign n37115 = n17629 & n37114;
  assign n37116 = n17765 & n37115;
  assign n37117 = n17874 & n37116;
  assign n37118 = ~n37108 & ~n37117;
  assign n37119 = n37096 & n37118;
  assign n37120 = n37072 & n37119;
  assign n37121 = n36989 & n37120;
  assign po136 = ~n36911 | ~n37121;
  assign n37123 = pi248 & ~n16144;
  assign n37124 = ~n16175 & n37123;
  assign n37125 = ~n16360 & n37124;
  assign n37126 = ~n17630 & n37125;
  assign n37127 = ~n16216 & n37126;
  assign n37128 = ~n16215 & n37127;
  assign n37129 = n16222 & n37128;
  assign n37130 = n17637 & n37129;
  assign n37131 = n17629 & n37130;
  assign n37132 = n17628 & n37131;
  assign n37133 = n17736 & n37132;
  assign n37134 = ~n780 & n26952;
  assign n37135 = ~n1372 & n37134;
  assign n37136 = ~n2243 & n37135;
  assign n37137 = ~n3104 & n37136;
  assign n37138 = ~n3971 & n37137;
  assign n37139 = ~n16682 & n37138;
  assign n37140 = ~n4872 & n37139;
  assign n37141 = ~n5801 & n37140;
  assign n37142 = ~n6739 & n37141;
  assign n37143 = ~n7807 & n37142;
  assign n37144 = ~n8989 & n37143;
  assign n37145 = ~n10273 & n37144;
  assign n37146 = ~n16680 & n37145;
  assign n37147 = ~n16679 & n37146;
  assign n37148 = ~n11499 & n37147;
  assign n37149 = ~n13076 & n37148;
  assign n37150 = ~n14698 & n37149;
  assign n37151 = ~n16678 & n37150;
  assign n37152 = ~n16677 & n37151;
  assign n37153 = n16704 & n37152;
  assign n37154 = n16707 & n37153;
  assign n37155 = n16711 & n37154;
  assign n37156 = n16676 & n37155;
  assign n37157 = n16736 & n37156;
  assign n37158 = ~n37133 & ~n37157;
  assign n37159 = ~n9763 & n34166;
  assign n37160 = ~n9929 & n37159;
  assign n37161 = ~n17263 & n37160;
  assign n37162 = ~n17262 & n37161;
  assign n37163 = ~n11266 & n37162;
  assign n37164 = ~n11588 & n37163;
  assign n37165 = ~n13859 & n37164;
  assign n37166 = ~n16216 & n37165;
  assign n37167 = ~n16215 & n37166;
  assign n37168 = n16222 & n37167;
  assign n37169 = n17273 & n37168;
  assign n37170 = n17277 & n37169;
  assign n37171 = n17261 & n37170;
  assign n37172 = n17302 & n37171;
  assign n37173 = pi216 & ~n12743;
  assign n37174 = ~n12773 & n37173;
  assign n37175 = ~n12902 & n37174;
  assign n37176 = ~n17419 & n37175;
  assign n37177 = ~n17418 & n37176;
  assign n37178 = ~n14009 & n37177;
  assign n37179 = ~n16216 & n37178;
  assign n37180 = ~n16215 & n37179;
  assign n37181 = n16222 & n37180;
  assign n37182 = n17427 & n37181;
  assign n37183 = n17431 & n37182;
  assign n37184 = n16214 & n37183;
  assign n37185 = n17456 & n37184;
  assign n37186 = ~n37172 & ~n37185;
  assign n37187 = n37158 & n37186;
  assign n37188 = ~n13820 & n34190;
  assign n37189 = ~n16216 & n37188;
  assign n37190 = ~n14741 & n37189;
  assign n37191 = ~n16209 & n37190;
  assign n37192 = ~n16211 & n37191;
  assign n37193 = n17238 & n37192;
  assign n37194 = n17232 & n37193;
  assign n37195 = n17225 & n37194;
  assign n37196 = ~n13906 & n34198;
  assign n37197 = ~n16216 & n37196;
  assign n37198 = ~n15586 & n37197;
  assign n37199 = ~n16208 & n37198;
  assign n37200 = n17257 & n37199;
  assign n37201 = n17328 & n37200;
  assign n37202 = n17342 & n37201;
  assign n37203 = ~n37195 & ~n37202;
  assign n37204 = ~n13093 & n31675;
  assign n37205 = ~n16216 & n37204;
  assign n37206 = ~n16215 & n37205;
  assign n37207 = n16222 & n37206;
  assign n37208 = n17516 & n37207;
  assign n37209 = n16214 & n37208;
  assign n37210 = n17512 & n37209;
  assign n37211 = n17534 & n37210;
  assign n37212 = ~n14073 & n34182;
  assign n37213 = ~n16216 & n37212;
  assign n37214 = ~n15616 & n37213;
  assign n37215 = ~n16224 & n37214;
  assign n37216 = n17086 & n37215;
  assign n37217 = n17351 & n37216;
  assign n37218 = n17350 & n37217;
  assign n37219 = n17370 & n37218;
  assign n37220 = ~n37211 & ~n37219;
  assign n37221 = n37203 & n37220;
  assign n37222 = ~n15075 & n34279;
  assign n37223 = ~n16216 & n37222;
  assign n37224 = ~n16537 & n37223;
  assign n37225 = n16544 & n37224;
  assign n37226 = ~n16831 & n34274;
  assign n37227 = ~n16829 & n37226;
  assign n37228 = n16836 & n37227;
  assign n37229 = pi264 & ~n501;
  assign n37230 = n12872 & n37229;
  assign n37231 = n17949 & n37230;
  assign n37232 = n17954 & n37231;
  assign n37233 = n17947 & n37232;
  assign n37234 = n17982 & n37233;
  assign n37235 = ~n1172 & n37234;
  assign n37236 = ~n996 & n37235;
  assign n37237 = ~n2306 & n37236;
  assign n37238 = ~n500 & n37237;
  assign n37239 = n17940 & n37238;
  assign n37240 = n17991 & n37239;
  assign n37241 = n17938 & n37240;
  assign n37242 = n17929 & n37241;
  assign n37243 = n17921 & n37242;
  assign n37244 = n18029 & n37243;
  assign n37245 = ~n7236 & n37244;
  assign n37246 = ~n6137 & n37245;
  assign n37247 = n6193 & n37246;
  assign n37248 = n6134 & n37247;
  assign n37249 = ~n8867 & n37248;
  assign n37250 = ~n7235 & n37249;
  assign n37251 = n7296 & n37250;
  assign n37252 = n7231 & n37251;
  assign n37253 = ~n10027 & n37252;
  assign n37254 = ~n8866 & n37253;
  assign n37255 = n8898 & n37254;
  assign n37256 = n8863 & n37255;
  assign n37257 = pi272 & ~n501;
  assign n37258 = n12872 & n37257;
  assign n37259 = n18049 & n37258;
  assign n37260 = n18053 & n37259;
  assign n37261 = n18047 & n37260;
  assign n37262 = n18080 & n37261;
  assign n37263 = ~n1172 & n37262;
  assign n37264 = ~n996 & n37263;
  assign n37265 = ~n2306 & n37264;
  assign n37266 = ~n500 & n37265;
  assign n37267 = n18038 & n37266;
  assign n37268 = n18037 & n37267;
  assign n37269 = n18088 & n37268;
  assign n37270 = n18106 & n37269;
  assign n37271 = n18035 & n37270;
  assign n37272 = n18134 & n37271;
  assign n37273 = ~n7236 & n37272;
  assign n37274 = ~n6137 & n37273;
  assign n37275 = n6193 & n37274;
  assign n37276 = n6134 & n37275;
  assign n37277 = ~n8867 & n37276;
  assign n37278 = ~n7235 & n37277;
  assign n37279 = n7296 & n37278;
  assign n37280 = n7231 & n37279;
  assign n37281 = ~n10027 & n37280;
  assign n37282 = ~n8866 & n37281;
  assign n37283 = n8898 & n37282;
  assign n37284 = n8863 & n37283;
  assign n37285 = ~n37256 & ~n37284;
  assign n37286 = ~n10788 & ~n37285;
  assign n37287 = ~n10026 & n37286;
  assign n37288 = n10072 & n37287;
  assign n37289 = n10021 & n37288;
  assign n37290 = ~n37228 & ~n37289;
  assign n37291 = ~n37225 & n37290;
  assign n37292 = ~n15278 & n34207;
  assign n37293 = ~n16216 & n37292;
  assign n37294 = n16939 & n37293;
  assign n37295 = ~n16937 & n37294;
  assign n37296 = n16944 & n37295;
  assign n37297 = n16936 & n37296;
  assign n37298 = ~n15167 & n34283;
  assign n37299 = ~n16216 & n37298;
  assign n37300 = ~n16220 & n37299;
  assign n37301 = ~n16466 & n37300;
  assign n37302 = n16476 & n37301;
  assign n37303 = ~n37297 & ~n37302;
  assign n37304 = n37291 & n37303;
  assign n37305 = ~n13764 & n34296;
  assign n37306 = ~n16216 & n37305;
  assign n37307 = ~n15465 & n37306;
  assign n37308 = ~n16209 & n37307;
  assign n37309 = n17086 & n37308;
  assign n37310 = n17133 & n37309;
  assign n37311 = n17122 & n37310;
  assign n37312 = ~n13726 & n34290;
  assign n37313 = ~n16216 & n37312;
  assign n37314 = ~n15419 & n37313;
  assign n37315 = n17086 & n37314;
  assign n37316 = n17094 & n37315;
  assign n37317 = n17083 & n37316;
  assign n37318 = ~n37311 & ~n37317;
  assign n37319 = n37304 & n37318;
  assign n37320 = n37221 & n37319;
  assign n37321 = n37187 & n37320;
  assign n37322 = pi120 & ~n5686;
  assign n37323 = ~n5349 & n37322;
  assign n37324 = ~n5808 & n37323;
  assign n37325 = ~n6056 & n37324;
  assign n37326 = ~n7073 & n37325;
  assign n37327 = ~n8179 & n37326;
  assign n37328 = ~n9344 & n37327;
  assign n37329 = ~n16418 & n37328;
  assign n37330 = ~n16361 & n37329;
  assign n37331 = ~n10594 & n37330;
  assign n37332 = ~n12005 & n37331;
  assign n37333 = ~n13558 & n37332;
  assign n37334 = ~n16216 & n37333;
  assign n37335 = ~n16215 & n37334;
  assign n37336 = n16432 & n37335;
  assign n37337 = n16435 & n37336;
  assign n37338 = n16439 & n37337;
  assign n37339 = n16305 & n37338;
  assign n37340 = n16464 & n37339;
  assign n37341 = pi072 & ~n2602;
  assign n37342 = ~n2783 & n37341;
  assign n37343 = ~n3066 & n37342;
  assign n37344 = ~n3983 & n37343;
  assign n37345 = ~n4003 & n37344;
  assign n37346 = ~n4024 & n37345;
  assign n37347 = ~n4999 & n37346;
  assign n37348 = ~n5827 & n37347;
  assign n37349 = ~n6893 & n37348;
  assign n37350 = ~n7890 & n37349;
  assign n37351 = ~n9131 & n37350;
  assign n37352 = ~n16617 & n37351;
  assign n37353 = ~n16616 & n37352;
  assign n37354 = ~n10278 & n37353;
  assign n37355 = ~n11662 & n37354;
  assign n37356 = ~n13191 & n37355;
  assign n37357 = ~n16615 & n37356;
  assign n37358 = ~n16614 & n37357;
  assign n37359 = n16636 & n37358;
  assign n37360 = n16639 & n37359;
  assign n37361 = n16643 & n37360;
  assign n37362 = n16613 & n37361;
  assign n37363 = n16668 & n37362;
  assign n37364 = ~n37340 & ~n37363;
  assign n37365 = pi168 & ~n8633;
  assign n37366 = ~n8455 & n37365;
  assign n37367 = ~n8834 & n37366;
  assign n37368 = ~n10002 & n37367;
  assign n37369 = ~n17152 & n37368;
  assign n37370 = ~n17151 & n37369;
  assign n37371 = ~n11297 & n37370;
  assign n37372 = ~n12240 & n37371;
  assign n37373 = ~n13135 & n37372;
  assign n37374 = ~n16216 & n37373;
  assign n37375 = ~n16215 & n37374;
  assign n37376 = n16222 & n37375;
  assign n37377 = n17163 & n37376;
  assign n37378 = n17167 & n37377;
  assign n37379 = n17150 & n37378;
  assign n37380 = n17192 & n37379;
  assign n37381 = ~n6401 & n27007;
  assign n37382 = ~n6784 & n37381;
  assign n37383 = ~n7158 & n37382;
  assign n37384 = ~n8250 & n37383;
  assign n37385 = ~n9414 & n37384;
  assign n37386 = ~n16957 & n37385;
  assign n37387 = ~n16956 & n37386;
  assign n37388 = ~n10667 & n37387;
  assign n37389 = ~n12083 & n37388;
  assign n37390 = ~n13644 & n37389;
  assign n37391 = ~n16216 & n37390;
  assign n37392 = ~n16215 & n37391;
  assign n37393 = n16222 & n37392;
  assign n37394 = n16971 & n37393;
  assign n37395 = n16975 & n37394;
  assign n37396 = n16955 & n37395;
  assign n37397 = n17000 & n37396;
  assign n37398 = ~n37380 & ~n37397;
  assign n37399 = n37364 & n37398;
  assign n37400 = pi256 & ~n16417;
  assign n37401 = ~n17766 & n37400;
  assign n37402 = ~n16216 & n37401;
  assign n37403 = ~n16215 & n37402;
  assign n37404 = n16222 & n37403;
  assign n37405 = n17637 & n37404;
  assign n37406 = n17629 & n37405;
  assign n37407 = n17765 & n37406;
  assign n37408 = n17874 & n37407;
  assign n37409 = ~n11042 & n34395;
  assign n37410 = ~n11188 & n37409;
  assign n37411 = ~n17378 & n37410;
  assign n37412 = ~n17377 & n37411;
  assign n37413 = ~n12380 & n37412;
  assign n37414 = ~n14045 & n37413;
  assign n37415 = ~n16216 & n37414;
  assign n37416 = ~n16215 & n37415;
  assign n37417 = n16222 & n37416;
  assign n37418 = n17387 & n37417;
  assign n37419 = n17391 & n37418;
  assign n37420 = n17376 & n37419;
  assign n37421 = n17416 & n37420;
  assign n37422 = ~n37408 & ~n37421;
  assign n37423 = ~n4460 & n34111;
  assign n37424 = ~n4817 & n37423;
  assign n37425 = ~n4902 & n37424;
  assign n37426 = ~n6001 & n37425;
  assign n37427 = ~n7014 & n37426;
  assign n37428 = ~n8114 & n37427;
  assign n37429 = ~n9276 & n37428;
  assign n37430 = ~n16486 & n37429;
  assign n37431 = ~n16485 & n37430;
  assign n37432 = ~n10523 & n37431;
  assign n37433 = ~n11928 & n37432;
  assign n37434 = ~n13479 & n37433;
  assign n37435 = ~n16216 & n37434;
  assign n37436 = ~n16220 & n37435;
  assign n37437 = n16503 & n37436;
  assign n37438 = n16506 & n37437;
  assign n37439 = n16510 & n37438;
  assign n37440 = n16484 & n37439;
  assign n37441 = n16535 & n37440;
  assign n37442 = pi056 & ~n1526;
  assign n37443 = ~n1556 & n37442;
  assign n37444 = ~n2242 & n37443;
  assign n37445 = ~n3095 & n37444;
  assign n37446 = ~n3997 & n37445;
  assign n37447 = ~n4003 & n37446;
  assign n37448 = ~n4837 & n37447;
  assign n37449 = ~n5822 & n37448;
  assign n37450 = ~n6820 & n37449;
  assign n37451 = ~n7785 & n37450;
  assign n37452 = ~n9027 & n37451;
  assign n37453 = ~n10245 & n37452;
  assign n37454 = ~n16748 & n37453;
  assign n37455 = ~n16747 & n37454;
  assign n37456 = ~n11536 & n37455;
  assign n37457 = ~n13036 & n37456;
  assign n37458 = ~n14653 & n37457;
  assign n37459 = ~n16746 & n37458;
  assign n37460 = ~n16745 & n37459;
  assign n37461 = n16770 & n37460;
  assign n37462 = n16773 & n37461;
  assign n37463 = n16777 & n37462;
  assign n37464 = n16744 & n37463;
  assign n37465 = n16802 & n37464;
  assign n37466 = ~n37441 & ~n37465;
  assign n37467 = n37422 & n37466;
  assign n37468 = ~n7505 & n23403;
  assign n37469 = ~n7869 & n37468;
  assign n37470 = ~n8346 & n37469;
  assign n37471 = ~n9485 & n37470;
  assign n37472 = ~n17018 & n37471;
  assign n37473 = ~n17017 & n37472;
  assign n37474 = ~n10741 & n37473;
  assign n37475 = ~n12158 & n37474;
  assign n37476 = ~n13693 & n37475;
  assign n37477 = ~n16216 & n37476;
  assign n37478 = ~n16215 & n37477;
  assign n37479 = n16222 & n37478;
  assign n37480 = n17031 & n37479;
  assign n37481 = n17035 & n37480;
  assign n37482 = n17016 & n37481;
  assign n37483 = n17060 & n37482;
  assign n37484 = ~n16216 & n34314;
  assign n37485 = ~n16215 & n37484;
  assign n37486 = n16222 & n37485;
  assign n37487 = n16225 & n37486;
  assign n37488 = n16229 & n37487;
  assign n37489 = n16214 & n37488;
  assign n37490 = n16297 & n37489;
  assign n37491 = ~n37483 & ~n37490;
  assign n37492 = ~n3650 & n26787;
  assign n37493 = ~n3940 & n37492;
  assign n37494 = ~n4001 & n37493;
  assign n37495 = ~n5043 & n37494;
  assign n37496 = ~n5943 & n37495;
  assign n37497 = ~n6951 & n37496;
  assign n37498 = ~n8037 & n37497;
  assign n37499 = ~n9200 & n37498;
  assign n37500 = ~n16555 & n37499;
  assign n37501 = ~n16554 & n37500;
  assign n37502 = ~n10445 & n37501;
  assign n37503 = ~n11846 & n37502;
  assign n37504 = ~n13393 & n37503;
  assign n37505 = ~n16216 & n37504;
  assign n37506 = ~n16553 & n37505;
  assign n37507 = n16573 & n37506;
  assign n37508 = n16576 & n37507;
  assign n37509 = n16580 & n37508;
  assign n37510 = n16552 & n37509;
  assign n37511 = n16605 & n37510;
  assign n37512 = pi232 & ~n14350;
  assign n37513 = ~n14381 & n37512;
  assign n37514 = ~n14519 & n37513;
  assign n37515 = ~n17537 & n37514;
  assign n37516 = ~n17536 & n37515;
  assign n37517 = ~n16216 & n37516;
  assign n37518 = ~n16215 & n37517;
  assign n37519 = n16222 & n37518;
  assign n37520 = n17544 & n37519;
  assign n37521 = n17547 & n37520;
  assign n37522 = n16214 & n37521;
  assign n37523 = n17572 & n37522;
  assign n37524 = ~n37511 & ~n37523;
  assign n37525 = n37491 & n37524;
  assign n37526 = n37467 & n37525;
  assign n37527 = n37399 & n37526;
  assign po137 = ~n37321 | ~n37527;
  assign n37529 = ~n3650 & n27270;
  assign n37530 = ~n3940 & n37529;
  assign n37531 = ~n4001 & n37530;
  assign n37532 = ~n5043 & n37531;
  assign n37533 = ~n5943 & n37532;
  assign n37534 = ~n6951 & n37533;
  assign n37535 = ~n8037 & n37534;
  assign n37536 = ~n9200 & n37535;
  assign n37537 = ~n16555 & n37536;
  assign n37538 = ~n16554 & n37537;
  assign n37539 = ~n10445 & n37538;
  assign n37540 = ~n11846 & n37539;
  assign n37541 = ~n13393 & n37540;
  assign n37542 = ~n16216 & n37541;
  assign n37543 = ~n16553 & n37542;
  assign n37544 = n16573 & n37543;
  assign n37545 = n16576 & n37544;
  assign n37546 = n16580 & n37545;
  assign n37547 = n16552 & n37546;
  assign n37548 = n16605 & n37547;
  assign n37549 = pi249 & ~n16144;
  assign n37550 = ~n16175 & n37549;
  assign n37551 = ~n16360 & n37550;
  assign n37552 = ~n17630 & n37551;
  assign n37553 = ~n16216 & n37552;
  assign n37554 = ~n16215 & n37553;
  assign n37555 = n16222 & n37554;
  assign n37556 = n17637 & n37555;
  assign n37557 = n17629 & n37556;
  assign n37558 = n17628 & n37557;
  assign n37559 = n17736 & n37558;
  assign n37560 = ~n37548 & ~n37559;
  assign n37561 = ~n780 & n27215;
  assign n37562 = ~n1372 & n37561;
  assign n37563 = ~n2243 & n37562;
  assign n37564 = ~n3104 & n37563;
  assign n37565 = ~n3971 & n37564;
  assign n37566 = ~n16682 & n37565;
  assign n37567 = ~n4872 & n37566;
  assign n37568 = ~n5801 & n37567;
  assign n37569 = ~n6739 & n37568;
  assign n37570 = ~n7807 & n37569;
  assign n37571 = ~n8989 & n37570;
  assign n37572 = ~n10273 & n37571;
  assign n37573 = ~n16680 & n37572;
  assign n37574 = ~n16679 & n37573;
  assign n37575 = ~n11499 & n37574;
  assign n37576 = ~n13076 & n37575;
  assign n37577 = ~n14698 & n37576;
  assign n37578 = ~n16678 & n37577;
  assign n37579 = ~n16677 & n37578;
  assign n37580 = n16704 & n37579;
  assign n37581 = n16707 & n37580;
  assign n37582 = n16711 & n37581;
  assign n37583 = n16676 & n37582;
  assign n37584 = n16736 & n37583;
  assign n37585 = pi217 & ~n12743;
  assign n37586 = ~n12773 & n37585;
  assign n37587 = ~n12902 & n37586;
  assign n37588 = ~n17419 & n37587;
  assign n37589 = ~n17418 & n37588;
  assign n37590 = ~n14009 & n37589;
  assign n37591 = ~n16216 & n37590;
  assign n37592 = ~n16215 & n37591;
  assign n37593 = n16222 & n37592;
  assign n37594 = n17427 & n37593;
  assign n37595 = n17431 & n37594;
  assign n37596 = n16214 & n37595;
  assign n37597 = n17456 & n37596;
  assign n37598 = ~n37584 & ~n37597;
  assign n37599 = n37560 & n37598;
  assign n37600 = ~n13906 & n34557;
  assign n37601 = ~n16216 & n37600;
  assign n37602 = ~n15586 & n37601;
  assign n37603 = ~n16208 & n37602;
  assign n37604 = n17257 & n37603;
  assign n37605 = n17328 & n37604;
  assign n37606 = n17342 & n37605;
  assign n37607 = ~n13820 & n34542;
  assign n37608 = ~n16216 & n37607;
  assign n37609 = ~n14741 & n37608;
  assign n37610 = ~n16209 & n37609;
  assign n37611 = ~n16211 & n37610;
  assign n37612 = n17238 & n37611;
  assign n37613 = n17232 & n37612;
  assign n37614 = n17225 & n37613;
  assign n37615 = ~n37606 & ~n37614;
  assign n37616 = ~n14073 & n34649;
  assign n37617 = ~n16216 & n37616;
  assign n37618 = ~n15616 & n37617;
  assign n37619 = ~n16224 & n37618;
  assign n37620 = n17086 & n37619;
  assign n37621 = n17351 & n37620;
  assign n37622 = n17350 & n37621;
  assign n37623 = n17370 & n37622;
  assign n37624 = ~n13093 & n32017;
  assign n37625 = ~n16216 & n37624;
  assign n37626 = ~n16215 & n37625;
  assign n37627 = n16222 & n37626;
  assign n37628 = n17516 & n37627;
  assign n37629 = n16214 & n37628;
  assign n37630 = n17512 & n37629;
  assign n37631 = n17534 & n37630;
  assign n37632 = ~n37623 & ~n37631;
  assign n37633 = n37615 & n37632;
  assign n37634 = ~n15075 & n34638;
  assign n37635 = ~n16216 & n37634;
  assign n37636 = ~n16537 & n37635;
  assign n37637 = n16544 & n37636;
  assign n37638 = ~n16831 & n34633;
  assign n37639 = ~n16829 & n37638;
  assign n37640 = n16836 & n37639;
  assign n37641 = pi265 & ~n501;
  assign n37642 = n12872 & n37641;
  assign n37643 = n17949 & n37642;
  assign n37644 = n17954 & n37643;
  assign n37645 = n17947 & n37644;
  assign n37646 = n17982 & n37645;
  assign n37647 = ~n1172 & n37646;
  assign n37648 = ~n996 & n37647;
  assign n37649 = ~n2306 & n37648;
  assign n37650 = ~n500 & n37649;
  assign n37651 = n17940 & n37650;
  assign n37652 = n17991 & n37651;
  assign n37653 = n17938 & n37652;
  assign n37654 = n17929 & n37653;
  assign n37655 = n17921 & n37654;
  assign n37656 = n18029 & n37655;
  assign n37657 = ~n7236 & n37656;
  assign n37658 = ~n6137 & n37657;
  assign n37659 = n6193 & n37658;
  assign n37660 = n6134 & n37659;
  assign n37661 = ~n8867 & n37660;
  assign n37662 = ~n7235 & n37661;
  assign n37663 = n7296 & n37662;
  assign n37664 = n7231 & n37663;
  assign n37665 = ~n10027 & n37664;
  assign n37666 = ~n8866 & n37665;
  assign n37667 = n8898 & n37666;
  assign n37668 = n8863 & n37667;
  assign n37669 = pi273 & ~n501;
  assign n37670 = n12872 & n37669;
  assign n37671 = n18049 & n37670;
  assign n37672 = n18053 & n37671;
  assign n37673 = n18047 & n37672;
  assign n37674 = n18080 & n37673;
  assign n37675 = ~n1172 & n37674;
  assign n37676 = ~n996 & n37675;
  assign n37677 = ~n2306 & n37676;
  assign n37678 = ~n500 & n37677;
  assign n37679 = n18038 & n37678;
  assign n37680 = n18037 & n37679;
  assign n37681 = n18088 & n37680;
  assign n37682 = n18106 & n37681;
  assign n37683 = n18035 & n37682;
  assign n37684 = n18134 & n37683;
  assign n37685 = ~n7236 & n37684;
  assign n37686 = ~n6137 & n37685;
  assign n37687 = n6193 & n37686;
  assign n37688 = n6134 & n37687;
  assign n37689 = ~n8867 & n37688;
  assign n37690 = ~n7235 & n37689;
  assign n37691 = n7296 & n37690;
  assign n37692 = n7231 & n37691;
  assign n37693 = ~n10027 & n37692;
  assign n37694 = ~n8866 & n37693;
  assign n37695 = n8898 & n37694;
  assign n37696 = n8863 & n37695;
  assign n37697 = ~n37668 & ~n37696;
  assign n37698 = ~n10788 & ~n37697;
  assign n37699 = ~n10026 & n37698;
  assign n37700 = n10072 & n37699;
  assign n37701 = n10021 & n37700;
  assign n37702 = ~n37640 & ~n37701;
  assign n37703 = ~n37637 & n37702;
  assign n37704 = ~n15278 & n34566;
  assign n37705 = ~n16216 & n37704;
  assign n37706 = n16939 & n37705;
  assign n37707 = ~n16937 & n37706;
  assign n37708 = n16944 & n37707;
  assign n37709 = n16936 & n37708;
  assign n37710 = ~n15167 & n34642;
  assign n37711 = ~n16216 & n37710;
  assign n37712 = ~n16220 & n37711;
  assign n37713 = ~n16466 & n37712;
  assign n37714 = n16476 & n37713;
  assign n37715 = ~n37709 & ~n37714;
  assign n37716 = n37703 & n37715;
  assign n37717 = ~n13764 & n34550;
  assign n37718 = ~n16216 & n37717;
  assign n37719 = ~n15465 & n37718;
  assign n37720 = ~n16209 & n37719;
  assign n37721 = n17086 & n37720;
  assign n37722 = n17133 & n37721;
  assign n37723 = n17122 & n37722;
  assign n37724 = ~n13726 & n34657;
  assign n37725 = ~n16216 & n37724;
  assign n37726 = ~n15419 & n37725;
  assign n37727 = n17086 & n37726;
  assign n37728 = n17094 & n37727;
  assign n37729 = n17083 & n37728;
  assign n37730 = ~n37723 & ~n37729;
  assign n37731 = n37716 & n37730;
  assign n37732 = n37633 & n37731;
  assign n37733 = n37599 & n37732;
  assign n37734 = pi057 & ~n1526;
  assign n37735 = ~n1556 & n37734;
  assign n37736 = ~n2242 & n37735;
  assign n37737 = ~n3095 & n37736;
  assign n37738 = ~n3997 & n37737;
  assign n37739 = ~n4003 & n37738;
  assign n37740 = ~n4837 & n37739;
  assign n37741 = ~n5822 & n37740;
  assign n37742 = ~n6820 & n37741;
  assign n37743 = ~n7785 & n37742;
  assign n37744 = ~n9027 & n37743;
  assign n37745 = ~n10245 & n37744;
  assign n37746 = ~n16748 & n37745;
  assign n37747 = ~n16747 & n37746;
  assign n37748 = ~n11536 & n37747;
  assign n37749 = ~n13036 & n37748;
  assign n37750 = ~n14653 & n37749;
  assign n37751 = ~n16746 & n37750;
  assign n37752 = ~n16745 & n37751;
  assign n37753 = n16770 & n37752;
  assign n37754 = n16773 & n37753;
  assign n37755 = n16777 & n37754;
  assign n37756 = n16744 & n37755;
  assign n37757 = n16802 & n37756;
  assign n37758 = pi169 & ~n8633;
  assign n37759 = ~n8455 & n37758;
  assign n37760 = ~n8834 & n37759;
  assign n37761 = ~n10002 & n37760;
  assign n37762 = ~n17152 & n37761;
  assign n37763 = ~n17151 & n37762;
  assign n37764 = ~n11297 & n37763;
  assign n37765 = ~n12240 & n37764;
  assign n37766 = ~n13135 & n37765;
  assign n37767 = ~n16216 & n37766;
  assign n37768 = ~n16215 & n37767;
  assign n37769 = n16222 & n37768;
  assign n37770 = n17163 & n37769;
  assign n37771 = n17167 & n37770;
  assign n37772 = n17150 & n37771;
  assign n37773 = n17192 & n37772;
  assign n37774 = ~n37757 & ~n37773;
  assign n37775 = ~n6401 & n27238;
  assign n37776 = ~n6784 & n37775;
  assign n37777 = ~n7158 & n37776;
  assign n37778 = ~n8250 & n37777;
  assign n37779 = ~n9414 & n37778;
  assign n37780 = ~n16957 & n37779;
  assign n37781 = ~n16956 & n37780;
  assign n37782 = ~n10667 & n37781;
  assign n37783 = ~n12083 & n37782;
  assign n37784 = ~n13644 & n37783;
  assign n37785 = ~n16216 & n37784;
  assign n37786 = ~n16215 & n37785;
  assign n37787 = n16222 & n37786;
  assign n37788 = n16971 & n37787;
  assign n37789 = n16975 & n37788;
  assign n37790 = n16955 & n37789;
  assign n37791 = n17000 & n37790;
  assign n37792 = ~n11042 & n34837;
  assign n37793 = ~n11188 & n37792;
  assign n37794 = ~n17378 & n37793;
  assign n37795 = ~n17377 & n37794;
  assign n37796 = ~n12380 & n37795;
  assign n37797 = ~n14045 & n37796;
  assign n37798 = ~n16216 & n37797;
  assign n37799 = ~n16215 & n37798;
  assign n37800 = n16222 & n37799;
  assign n37801 = n17387 & n37800;
  assign n37802 = n17391 & n37801;
  assign n37803 = n17376 & n37802;
  assign n37804 = n17416 & n37803;
  assign n37805 = ~n37791 & ~n37804;
  assign n37806 = n37774 & n37805;
  assign n37807 = pi233 & ~n14350;
  assign n37808 = ~n14381 & n37807;
  assign n37809 = ~n14519 & n37808;
  assign n37810 = ~n17537 & n37809;
  assign n37811 = ~n17536 & n37810;
  assign n37812 = ~n16216 & n37811;
  assign n37813 = ~n16215 & n37812;
  assign n37814 = n16222 & n37813;
  assign n37815 = n17544 & n37814;
  assign n37816 = n17547 & n37815;
  assign n37817 = n16214 & n37816;
  assign n37818 = n17572 & n37817;
  assign n37819 = ~n9763 & n34704;
  assign n37820 = ~n9929 & n37819;
  assign n37821 = ~n17263 & n37820;
  assign n37822 = ~n17262 & n37821;
  assign n37823 = ~n11266 & n37822;
  assign n37824 = ~n11588 & n37823;
  assign n37825 = ~n13859 & n37824;
  assign n37826 = ~n16216 & n37825;
  assign n37827 = ~n16215 & n37826;
  assign n37828 = n16222 & n37827;
  assign n37829 = n17273 & n37828;
  assign n37830 = n17277 & n37829;
  assign n37831 = n17261 & n37830;
  assign n37832 = n17302 & n37831;
  assign n37833 = ~n37818 & ~n37832;
  assign n37834 = pi121 & ~n5686;
  assign n37835 = ~n5349 & n37834;
  assign n37836 = ~n5808 & n37835;
  assign n37837 = ~n6056 & n37836;
  assign n37838 = ~n7073 & n37837;
  assign n37839 = ~n8179 & n37838;
  assign n37840 = ~n9344 & n37839;
  assign n37841 = ~n16418 & n37840;
  assign n37842 = ~n16361 & n37841;
  assign n37843 = ~n10594 & n37842;
  assign n37844 = ~n12005 & n37843;
  assign n37845 = ~n13558 & n37844;
  assign n37846 = ~n16216 & n37845;
  assign n37847 = ~n16215 & n37846;
  assign n37848 = n16432 & n37847;
  assign n37849 = n16435 & n37848;
  assign n37850 = n16439 & n37849;
  assign n37851 = n16305 & n37850;
  assign n37852 = n16464 & n37851;
  assign n37853 = ~n4460 & n34720;
  assign n37854 = ~n4817 & n37853;
  assign n37855 = ~n4902 & n37854;
  assign n37856 = ~n6001 & n37855;
  assign n37857 = ~n7014 & n37856;
  assign n37858 = ~n8114 & n37857;
  assign n37859 = ~n9276 & n37858;
  assign n37860 = ~n16486 & n37859;
  assign n37861 = ~n16485 & n37860;
  assign n37862 = ~n10523 & n37861;
  assign n37863 = ~n11928 & n37862;
  assign n37864 = ~n13479 & n37863;
  assign n37865 = ~n16216 & n37864;
  assign n37866 = ~n16220 & n37865;
  assign n37867 = n16503 & n37866;
  assign n37868 = n16506 & n37867;
  assign n37869 = n16510 & n37868;
  assign n37870 = n16484 & n37869;
  assign n37871 = n16535 & n37870;
  assign n37872 = ~n37852 & ~n37871;
  assign n37873 = n37833 & n37872;
  assign n37874 = ~n7505 & n23526;
  assign n37875 = ~n7869 & n37874;
  assign n37876 = ~n8346 & n37875;
  assign n37877 = ~n9485 & n37876;
  assign n37878 = ~n17018 & n37877;
  assign n37879 = ~n17017 & n37878;
  assign n37880 = ~n10741 & n37879;
  assign n37881 = ~n12158 & n37880;
  assign n37882 = ~n13693 & n37881;
  assign n37883 = ~n16216 & n37882;
  assign n37884 = ~n16215 & n37883;
  assign n37885 = n16222 & n37884;
  assign n37886 = n17031 & n37885;
  assign n37887 = n17035 & n37886;
  assign n37888 = n17016 & n37887;
  assign n37889 = n17060 & n37888;
  assign n37890 = ~n16216 & n34770;
  assign n37891 = ~n16215 & n37890;
  assign n37892 = n16222 & n37891;
  assign n37893 = n16225 & n37892;
  assign n37894 = n16229 & n37893;
  assign n37895 = n16214 & n37894;
  assign n37896 = n16297 & n37895;
  assign n37897 = ~n37889 & ~n37896;
  assign n37898 = pi257 & ~n16417;
  assign n37899 = ~n17766 & n37898;
  assign n37900 = ~n16216 & n37899;
  assign n37901 = ~n16215 & n37900;
  assign n37902 = n16222 & n37901;
  assign n37903 = n17637 & n37902;
  assign n37904 = n17629 & n37903;
  assign n37905 = n17765 & n37904;
  assign n37906 = n17874 & n37905;
  assign n37907 = pi073 & ~n2602;
  assign n37908 = ~n2783 & n37907;
  assign n37909 = ~n3066 & n37908;
  assign n37910 = ~n3983 & n37909;
  assign n37911 = ~n4003 & n37910;
  assign n37912 = ~n4024 & n37911;
  assign n37913 = ~n4999 & n37912;
  assign n37914 = ~n5827 & n37913;
  assign n37915 = ~n6893 & n37914;
  assign n37916 = ~n7890 & n37915;
  assign n37917 = ~n9131 & n37916;
  assign n37918 = ~n16617 & n37917;
  assign n37919 = ~n16616 & n37918;
  assign n37920 = ~n10278 & n37919;
  assign n37921 = ~n11662 & n37920;
  assign n37922 = ~n13191 & n37921;
  assign n37923 = ~n16615 & n37922;
  assign n37924 = ~n16614 & n37923;
  assign n37925 = n16636 & n37924;
  assign n37926 = n16639 & n37925;
  assign n37927 = n16643 & n37926;
  assign n37928 = n16613 & n37927;
  assign n37929 = n16668 & n37928;
  assign n37930 = ~n37906 & ~n37929;
  assign n37931 = n37897 & n37930;
  assign n37932 = n37873 & n37931;
  assign n37933 = n37806 & n37932;
  assign po138 = ~n37733 | ~n37933;
  assign n37935 = ~n3650 & n27506;
  assign n37936 = ~n3940 & n37935;
  assign n37937 = ~n4001 & n37936;
  assign n37938 = ~n5043 & n37937;
  assign n37939 = ~n5943 & n37938;
  assign n37940 = ~n6951 & n37939;
  assign n37941 = ~n8037 & n37940;
  assign n37942 = ~n9200 & n37941;
  assign n37943 = ~n16555 & n37942;
  assign n37944 = ~n16554 & n37943;
  assign n37945 = ~n10445 & n37944;
  assign n37946 = ~n11846 & n37945;
  assign n37947 = ~n13393 & n37946;
  assign n37948 = ~n16216 & n37947;
  assign n37949 = ~n16553 & n37948;
  assign n37950 = n16573 & n37949;
  assign n37951 = n16576 & n37950;
  assign n37952 = n16580 & n37951;
  assign n37953 = n16552 & n37952;
  assign n37954 = n16605 & n37953;
  assign n37955 = pi250 & ~n16144;
  assign n37956 = ~n16175 & n37955;
  assign n37957 = ~n16360 & n37956;
  assign n37958 = ~n17630 & n37957;
  assign n37959 = ~n16216 & n37958;
  assign n37960 = ~n16215 & n37959;
  assign n37961 = n16222 & n37960;
  assign n37962 = n17637 & n37961;
  assign n37963 = n17629 & n37962;
  assign n37964 = n17628 & n37963;
  assign n37965 = n17736 & n37964;
  assign n37966 = ~n37954 & ~n37965;
  assign n37967 = ~n780 & n27477;
  assign n37968 = ~n1372 & n37967;
  assign n37969 = ~n2243 & n37968;
  assign n37970 = ~n3104 & n37969;
  assign n37971 = ~n3971 & n37970;
  assign n37972 = ~n16682 & n37971;
  assign n37973 = ~n4872 & n37972;
  assign n37974 = ~n5801 & n37973;
  assign n37975 = ~n6739 & n37974;
  assign n37976 = ~n7807 & n37975;
  assign n37977 = ~n8989 & n37976;
  assign n37978 = ~n10273 & n37977;
  assign n37979 = ~n16680 & n37978;
  assign n37980 = ~n16679 & n37979;
  assign n37981 = ~n11499 & n37980;
  assign n37982 = ~n13076 & n37981;
  assign n37983 = ~n14698 & n37982;
  assign n37984 = ~n16678 & n37983;
  assign n37985 = ~n16677 & n37984;
  assign n37986 = n16704 & n37985;
  assign n37987 = n16707 & n37986;
  assign n37988 = n16711 & n37987;
  assign n37989 = n16676 & n37988;
  assign n37990 = n16736 & n37989;
  assign n37991 = pi218 & ~n12743;
  assign n37992 = ~n12773 & n37991;
  assign n37993 = ~n12902 & n37992;
  assign n37994 = ~n17419 & n37993;
  assign n37995 = ~n17418 & n37994;
  assign n37996 = ~n14009 & n37995;
  assign n37997 = ~n16216 & n37996;
  assign n37998 = ~n16215 & n37997;
  assign n37999 = n16222 & n37998;
  assign n38000 = n17427 & n37999;
  assign n38001 = n17431 & n38000;
  assign n38002 = n16214 & n38001;
  assign n38003 = n17456 & n38002;
  assign n38004 = ~n37990 & ~n38003;
  assign n38005 = n37966 & n38004;
  assign n38006 = ~n13906 & n34923;
  assign n38007 = ~n16216 & n38006;
  assign n38008 = ~n15586 & n38007;
  assign n38009 = ~n16208 & n38008;
  assign n38010 = n17257 & n38009;
  assign n38011 = n17328 & n38010;
  assign n38012 = n17342 & n38011;
  assign n38013 = ~n13820 & n34915;
  assign n38014 = ~n16216 & n38013;
  assign n38015 = ~n14741 & n38014;
  assign n38016 = ~n16209 & n38015;
  assign n38017 = ~n16211 & n38016;
  assign n38018 = n17238 & n38017;
  assign n38019 = n17232 & n38018;
  assign n38020 = n17225 & n38019;
  assign n38021 = ~n38012 & ~n38020;
  assign n38022 = ~n14073 & n34930;
  assign n38023 = ~n16216 & n38022;
  assign n38024 = ~n15616 & n38023;
  assign n38025 = ~n16224 & n38024;
  assign n38026 = n17086 & n38025;
  assign n38027 = n17351 & n38026;
  assign n38028 = n17350 & n38027;
  assign n38029 = n17370 & n38028;
  assign n38030 = ~n13093 & n32388;
  assign n38031 = ~n16216 & n38030;
  assign n38032 = ~n16215 & n38031;
  assign n38033 = n16222 & n38032;
  assign n38034 = n17516 & n38033;
  assign n38035 = n16214 & n38034;
  assign n38036 = n17512 & n38035;
  assign n38037 = n17534 & n38036;
  assign n38038 = ~n38029 & ~n38037;
  assign n38039 = n38021 & n38038;
  assign n38040 = ~n15075 & n35012;
  assign n38041 = ~n16216 & n38040;
  assign n38042 = ~n16537 & n38041;
  assign n38043 = n16544 & n38042;
  assign n38044 = ~n16831 & n35007;
  assign n38045 = ~n16829 & n38044;
  assign n38046 = n16836 & n38045;
  assign n38047 = pi266 & ~n501;
  assign n38048 = n12872 & n38047;
  assign n38049 = n17949 & n38048;
  assign n38050 = n17954 & n38049;
  assign n38051 = n17947 & n38050;
  assign n38052 = n17982 & n38051;
  assign n38053 = ~n1172 & n38052;
  assign n38054 = ~n996 & n38053;
  assign n38055 = ~n2306 & n38054;
  assign n38056 = ~n500 & n38055;
  assign n38057 = n17940 & n38056;
  assign n38058 = n17991 & n38057;
  assign n38059 = n17938 & n38058;
  assign n38060 = n17929 & n38059;
  assign n38061 = n17921 & n38060;
  assign n38062 = n18029 & n38061;
  assign n38063 = ~n7236 & n38062;
  assign n38064 = ~n6137 & n38063;
  assign n38065 = n6193 & n38064;
  assign n38066 = n6134 & n38065;
  assign n38067 = ~n8867 & n38066;
  assign n38068 = ~n7235 & n38067;
  assign n38069 = n7296 & n38068;
  assign n38070 = n7231 & n38069;
  assign n38071 = ~n10027 & n38070;
  assign n38072 = ~n8866 & n38071;
  assign n38073 = n8898 & n38072;
  assign n38074 = n8863 & n38073;
  assign n38075 = pi274 & ~n501;
  assign n38076 = n12872 & n38075;
  assign n38077 = n18049 & n38076;
  assign n38078 = n18053 & n38077;
  assign n38079 = n18047 & n38078;
  assign n38080 = n18080 & n38079;
  assign n38081 = ~n1172 & n38080;
  assign n38082 = ~n996 & n38081;
  assign n38083 = ~n2306 & n38082;
  assign n38084 = ~n500 & n38083;
  assign n38085 = n18038 & n38084;
  assign n38086 = n18037 & n38085;
  assign n38087 = n18088 & n38086;
  assign n38088 = n18106 & n38087;
  assign n38089 = n18035 & n38088;
  assign n38090 = n18134 & n38089;
  assign n38091 = ~n7236 & n38090;
  assign n38092 = ~n6137 & n38091;
  assign n38093 = n6193 & n38092;
  assign n38094 = n6134 & n38093;
  assign n38095 = ~n8867 & n38094;
  assign n38096 = ~n7235 & n38095;
  assign n38097 = n7296 & n38096;
  assign n38098 = n7231 & n38097;
  assign n38099 = ~n10027 & n38098;
  assign n38100 = ~n8866 & n38099;
  assign n38101 = n8898 & n38100;
  assign n38102 = n8863 & n38101;
  assign n38103 = ~n38074 & ~n38102;
  assign n38104 = ~n10788 & ~n38103;
  assign n38105 = ~n10026 & n38104;
  assign n38106 = n10072 & n38105;
  assign n38107 = n10021 & n38106;
  assign n38108 = ~n38046 & ~n38107;
  assign n38109 = ~n38043 & n38108;
  assign n38110 = ~n15278 & n34940;
  assign n38111 = ~n16216 & n38110;
  assign n38112 = n16939 & n38111;
  assign n38113 = ~n16937 & n38112;
  assign n38114 = n16944 & n38113;
  assign n38115 = n16936 & n38114;
  assign n38116 = ~n15167 & n35016;
  assign n38117 = ~n16216 & n38116;
  assign n38118 = ~n16220 & n38117;
  assign n38119 = ~n16466 & n38118;
  assign n38120 = n16476 & n38119;
  assign n38121 = ~n38115 & ~n38120;
  assign n38122 = n38109 & n38121;
  assign n38123 = ~n13764 & n35023;
  assign n38124 = ~n16216 & n38123;
  assign n38125 = ~n15465 & n38124;
  assign n38126 = ~n16209 & n38125;
  assign n38127 = n17086 & n38126;
  assign n38128 = n17133 & n38127;
  assign n38129 = n17122 & n38128;
  assign n38130 = ~n13726 & n35030;
  assign n38131 = ~n16216 & n38130;
  assign n38132 = ~n15419 & n38131;
  assign n38133 = n17086 & n38132;
  assign n38134 = n17094 & n38133;
  assign n38135 = n17083 & n38134;
  assign n38136 = ~n38129 & ~n38135;
  assign n38137 = n38122 & n38136;
  assign n38138 = n38039 & n38137;
  assign n38139 = n38005 & n38138;
  assign n38140 = pi258 & ~n16417;
  assign n38141 = ~n17766 & n38140;
  assign n38142 = ~n16216 & n38141;
  assign n38143 = ~n16215 & n38142;
  assign n38144 = n16222 & n38143;
  assign n38145 = n17637 & n38144;
  assign n38146 = n17629 & n38145;
  assign n38147 = n17765 & n38146;
  assign n38148 = n17874 & n38147;
  assign n38149 = pi170 & ~n8633;
  assign n38150 = ~n8455 & n38149;
  assign n38151 = ~n8834 & n38150;
  assign n38152 = ~n10002 & n38151;
  assign n38153 = ~n17152 & n38152;
  assign n38154 = ~n17151 & n38153;
  assign n38155 = ~n11297 & n38154;
  assign n38156 = ~n12240 & n38155;
  assign n38157 = ~n13135 & n38156;
  assign n38158 = ~n16216 & n38157;
  assign n38159 = ~n16215 & n38158;
  assign n38160 = n16222 & n38159;
  assign n38161 = n17163 & n38160;
  assign n38162 = n17167 & n38161;
  assign n38163 = n17150 & n38162;
  assign n38164 = n17192 & n38163;
  assign n38165 = ~n38148 & ~n38164;
  assign n38166 = ~n6401 & n27435;
  assign n38167 = ~n6784 & n38166;
  assign n38168 = ~n7158 & n38167;
  assign n38169 = ~n8250 & n38168;
  assign n38170 = ~n9414 & n38169;
  assign n38171 = ~n16957 & n38170;
  assign n38172 = ~n16956 & n38171;
  assign n38173 = ~n10667 & n38172;
  assign n38174 = ~n12083 & n38173;
  assign n38175 = ~n13644 & n38174;
  assign n38176 = ~n16216 & n38175;
  assign n38177 = ~n16215 & n38176;
  assign n38178 = n16222 & n38177;
  assign n38179 = n16971 & n38178;
  assign n38180 = n16975 & n38179;
  assign n38181 = n16955 & n38180;
  assign n38182 = n17000 & n38181;
  assign n38183 = ~n11042 & n35197;
  assign n38184 = ~n11188 & n38183;
  assign n38185 = ~n17378 & n38184;
  assign n38186 = ~n17377 & n38185;
  assign n38187 = ~n12380 & n38186;
  assign n38188 = ~n14045 & n38187;
  assign n38189 = ~n16216 & n38188;
  assign n38190 = ~n16215 & n38189;
  assign n38191 = n16222 & n38190;
  assign n38192 = n17387 & n38191;
  assign n38193 = n17391 & n38192;
  assign n38194 = n17376 & n38193;
  assign n38195 = n17416 & n38194;
  assign n38196 = ~n38182 & ~n38195;
  assign n38197 = n38165 & n38196;
  assign n38198 = ~n9763 & n35077;
  assign n38199 = ~n9929 & n38198;
  assign n38200 = ~n17263 & n38199;
  assign n38201 = ~n17262 & n38200;
  assign n38202 = ~n11266 & n38201;
  assign n38203 = ~n11588 & n38202;
  assign n38204 = ~n13859 & n38203;
  assign n38205 = ~n16216 & n38204;
  assign n38206 = ~n16215 & n38205;
  assign n38207 = n16222 & n38206;
  assign n38208 = n17273 & n38207;
  assign n38209 = n17277 & n38208;
  assign n38210 = n17261 & n38209;
  assign n38211 = n17302 & n38210;
  assign n38212 = pi122 & ~n5686;
  assign n38213 = ~n5349 & n38212;
  assign n38214 = ~n5808 & n38213;
  assign n38215 = ~n6056 & n38214;
  assign n38216 = ~n7073 & n38215;
  assign n38217 = ~n8179 & n38216;
  assign n38218 = ~n9344 & n38217;
  assign n38219 = ~n16418 & n38218;
  assign n38220 = ~n16361 & n38219;
  assign n38221 = ~n10594 & n38220;
  assign n38222 = ~n12005 & n38221;
  assign n38223 = ~n13558 & n38222;
  assign n38224 = ~n16216 & n38223;
  assign n38225 = ~n16215 & n38224;
  assign n38226 = n16432 & n38225;
  assign n38227 = n16435 & n38226;
  assign n38228 = n16439 & n38227;
  assign n38229 = n16305 & n38228;
  assign n38230 = n16464 & n38229;
  assign n38231 = ~n38211 & ~n38230;
  assign n38232 = ~n4460 & n35128;
  assign n38233 = ~n4817 & n38232;
  assign n38234 = ~n4902 & n38233;
  assign n38235 = ~n6001 & n38234;
  assign n38236 = ~n7014 & n38235;
  assign n38237 = ~n8114 & n38236;
  assign n38238 = ~n9276 & n38237;
  assign n38239 = ~n16486 & n38238;
  assign n38240 = ~n16485 & n38239;
  assign n38241 = ~n10523 & n38240;
  assign n38242 = ~n11928 & n38241;
  assign n38243 = ~n13479 & n38242;
  assign n38244 = ~n16216 & n38243;
  assign n38245 = ~n16220 & n38244;
  assign n38246 = n16503 & n38245;
  assign n38247 = n16506 & n38246;
  assign n38248 = n16510 & n38247;
  assign n38249 = n16484 & n38248;
  assign n38250 = n16535 & n38249;
  assign n38251 = pi058 & ~n1526;
  assign n38252 = ~n1556 & n38251;
  assign n38253 = ~n2242 & n38252;
  assign n38254 = ~n3095 & n38253;
  assign n38255 = ~n3997 & n38254;
  assign n38256 = ~n4003 & n38255;
  assign n38257 = ~n4837 & n38256;
  assign n38258 = ~n5822 & n38257;
  assign n38259 = ~n6820 & n38258;
  assign n38260 = ~n7785 & n38259;
  assign n38261 = ~n9027 & n38260;
  assign n38262 = ~n10245 & n38261;
  assign n38263 = ~n16748 & n38262;
  assign n38264 = ~n16747 & n38263;
  assign n38265 = ~n11536 & n38264;
  assign n38266 = ~n13036 & n38265;
  assign n38267 = ~n14653 & n38266;
  assign n38268 = ~n16746 & n38267;
  assign n38269 = ~n16745 & n38268;
  assign n38270 = n16770 & n38269;
  assign n38271 = n16773 & n38270;
  assign n38272 = n16777 & n38271;
  assign n38273 = n16744 & n38272;
  assign n38274 = n16802 & n38273;
  assign n38275 = ~n38250 & ~n38274;
  assign n38276 = n38231 & n38275;
  assign n38277 = ~n7505 & n23752;
  assign n38278 = ~n7869 & n38277;
  assign n38279 = ~n8346 & n38278;
  assign n38280 = ~n9485 & n38279;
  assign n38281 = ~n17018 & n38280;
  assign n38282 = ~n17017 & n38281;
  assign n38283 = ~n10741 & n38282;
  assign n38284 = ~n12158 & n38283;
  assign n38285 = ~n13693 & n38284;
  assign n38286 = ~n16216 & n38285;
  assign n38287 = ~n16215 & n38286;
  assign n38288 = n16222 & n38287;
  assign n38289 = n17031 & n38288;
  assign n38290 = n17035 & n38289;
  assign n38291 = n17016 & n38290;
  assign n38292 = n17060 & n38291;
  assign n38293 = ~n16216 & n35172;
  assign n38294 = ~n16215 & n38293;
  assign n38295 = n16222 & n38294;
  assign n38296 = n16225 & n38295;
  assign n38297 = n16229 & n38296;
  assign n38298 = n16214 & n38297;
  assign n38299 = n16297 & n38298;
  assign n38300 = ~n38292 & ~n38299;
  assign n38301 = pi074 & ~n2602;
  assign n38302 = ~n2783 & n38301;
  assign n38303 = ~n3066 & n38302;
  assign n38304 = ~n3983 & n38303;
  assign n38305 = ~n4003 & n38304;
  assign n38306 = ~n4024 & n38305;
  assign n38307 = ~n4999 & n38306;
  assign n38308 = ~n5827 & n38307;
  assign n38309 = ~n6893 & n38308;
  assign n38310 = ~n7890 & n38309;
  assign n38311 = ~n9131 & n38310;
  assign n38312 = ~n16617 & n38311;
  assign n38313 = ~n16616 & n38312;
  assign n38314 = ~n10278 & n38313;
  assign n38315 = ~n11662 & n38314;
  assign n38316 = ~n13191 & n38315;
  assign n38317 = ~n16615 & n38316;
  assign n38318 = ~n16614 & n38317;
  assign n38319 = n16636 & n38318;
  assign n38320 = n16639 & n38319;
  assign n38321 = n16643 & n38320;
  assign n38322 = n16613 & n38321;
  assign n38323 = n16668 & n38322;
  assign n38324 = pi234 & ~n14350;
  assign n38325 = ~n14381 & n38324;
  assign n38326 = ~n14519 & n38325;
  assign n38327 = ~n17537 & n38326;
  assign n38328 = ~n17536 & n38327;
  assign n38329 = ~n16216 & n38328;
  assign n38330 = ~n16215 & n38329;
  assign n38331 = n16222 & n38330;
  assign n38332 = n17544 & n38331;
  assign n38333 = n17547 & n38332;
  assign n38334 = n16214 & n38333;
  assign n38335 = n17572 & n38334;
  assign n38336 = ~n38323 & ~n38335;
  assign n38337 = n38300 & n38336;
  assign n38338 = n38276 & n38337;
  assign n38339 = n38197 & n38338;
  assign po139 = ~n38139 | ~n38339;
  assign n38341 = ~n3650 & n27770;
  assign n38342 = ~n3940 & n38341;
  assign n38343 = ~n4001 & n38342;
  assign n38344 = ~n5043 & n38343;
  assign n38345 = ~n5943 & n38344;
  assign n38346 = ~n6951 & n38345;
  assign n38347 = ~n8037 & n38346;
  assign n38348 = ~n9200 & n38347;
  assign n38349 = ~n16555 & n38348;
  assign n38350 = ~n16554 & n38349;
  assign n38351 = ~n10445 & n38350;
  assign n38352 = ~n11846 & n38351;
  assign n38353 = ~n13393 & n38352;
  assign n38354 = ~n16216 & n38353;
  assign n38355 = ~n16553 & n38354;
  assign n38356 = n16573 & n38355;
  assign n38357 = n16576 & n38356;
  assign n38358 = n16580 & n38357;
  assign n38359 = n16552 & n38358;
  assign n38360 = n16605 & n38359;
  assign n38361 = pi251 & ~n16144;
  assign n38362 = ~n16175 & n38361;
  assign n38363 = ~n16360 & n38362;
  assign n38364 = ~n17630 & n38363;
  assign n38365 = ~n16216 & n38364;
  assign n38366 = ~n16215 & n38365;
  assign n38367 = n16222 & n38366;
  assign n38368 = n17637 & n38367;
  assign n38369 = n17629 & n38368;
  assign n38370 = n17628 & n38369;
  assign n38371 = n17736 & n38370;
  assign n38372 = ~n38360 & ~n38371;
  assign n38373 = ~n780 & n27731;
  assign n38374 = ~n1372 & n38373;
  assign n38375 = ~n2243 & n38374;
  assign n38376 = ~n3104 & n38375;
  assign n38377 = ~n3971 & n38376;
  assign n38378 = ~n16682 & n38377;
  assign n38379 = ~n4872 & n38378;
  assign n38380 = ~n5801 & n38379;
  assign n38381 = ~n6739 & n38380;
  assign n38382 = ~n7807 & n38381;
  assign n38383 = ~n8989 & n38382;
  assign n38384 = ~n10273 & n38383;
  assign n38385 = ~n16680 & n38384;
  assign n38386 = ~n16679 & n38385;
  assign n38387 = ~n11499 & n38386;
  assign n38388 = ~n13076 & n38387;
  assign n38389 = ~n14698 & n38388;
  assign n38390 = ~n16678 & n38389;
  assign n38391 = ~n16677 & n38390;
  assign n38392 = n16704 & n38391;
  assign n38393 = n16707 & n38392;
  assign n38394 = n16711 & n38393;
  assign n38395 = n16676 & n38394;
  assign n38396 = n16736 & n38395;
  assign n38397 = pi219 & ~n12743;
  assign n38398 = ~n12773 & n38397;
  assign n38399 = ~n12902 & n38398;
  assign n38400 = ~n17419 & n38399;
  assign n38401 = ~n17418 & n38400;
  assign n38402 = ~n14009 & n38401;
  assign n38403 = ~n16216 & n38402;
  assign n38404 = ~n16215 & n38403;
  assign n38405 = n16222 & n38404;
  assign n38406 = n17427 & n38405;
  assign n38407 = n17431 & n38406;
  assign n38408 = n16214 & n38407;
  assign n38409 = n17456 & n38408;
  assign n38410 = ~n38396 & ~n38409;
  assign n38411 = n38372 & n38410;
  assign n38412 = ~n13906 & n35307;
  assign n38413 = ~n16216 & n38412;
  assign n38414 = ~n15586 & n38413;
  assign n38415 = ~n16208 & n38414;
  assign n38416 = n17257 & n38415;
  assign n38417 = n17328 & n38416;
  assign n38418 = n17342 & n38417;
  assign n38419 = ~n13820 & n35299;
  assign n38420 = ~n16216 & n38419;
  assign n38421 = ~n14741 & n38420;
  assign n38422 = ~n16209 & n38421;
  assign n38423 = ~n16211 & n38422;
  assign n38424 = n17238 & n38423;
  assign n38425 = n17232 & n38424;
  assign n38426 = n17225 & n38425;
  assign n38427 = ~n38418 & ~n38426;
  assign n38428 = ~n14073 & n35399;
  assign n38429 = ~n16216 & n38428;
  assign n38430 = ~n15616 & n38429;
  assign n38431 = ~n16224 & n38430;
  assign n38432 = n17086 & n38431;
  assign n38433 = n17351 & n38432;
  assign n38434 = n17350 & n38433;
  assign n38435 = n17370 & n38434;
  assign n38436 = ~n13093 & n32576;
  assign n38437 = ~n16216 & n38436;
  assign n38438 = ~n16215 & n38437;
  assign n38439 = n16222 & n38438;
  assign n38440 = n17516 & n38439;
  assign n38441 = n16214 & n38440;
  assign n38442 = n17512 & n38441;
  assign n38443 = n17534 & n38442;
  assign n38444 = ~n38435 & ~n38443;
  assign n38445 = n38427 & n38444;
  assign n38446 = ~n15075 & n35316;
  assign n38447 = ~n16216 & n38446;
  assign n38448 = ~n16537 & n38447;
  assign n38449 = n16544 & n38448;
  assign n38450 = ~n16831 & n35320;
  assign n38451 = ~n16829 & n38450;
  assign n38452 = n16836 & n38451;
  assign n38453 = pi267 & ~n501;
  assign n38454 = n12872 & n38453;
  assign n38455 = n17949 & n38454;
  assign n38456 = n17954 & n38455;
  assign n38457 = n17947 & n38456;
  assign n38458 = n17982 & n38457;
  assign n38459 = ~n1172 & n38458;
  assign n38460 = ~n996 & n38459;
  assign n38461 = ~n2306 & n38460;
  assign n38462 = ~n500 & n38461;
  assign n38463 = n17940 & n38462;
  assign n38464 = n17991 & n38463;
  assign n38465 = n17938 & n38464;
  assign n38466 = n17929 & n38465;
  assign n38467 = n17921 & n38466;
  assign n38468 = n18029 & n38467;
  assign n38469 = ~n7236 & n38468;
  assign n38470 = ~n6137 & n38469;
  assign n38471 = n6193 & n38470;
  assign n38472 = n6134 & n38471;
  assign n38473 = ~n8867 & n38472;
  assign n38474 = ~n7235 & n38473;
  assign n38475 = n7296 & n38474;
  assign n38476 = n7231 & n38475;
  assign n38477 = ~n10027 & n38476;
  assign n38478 = ~n8866 & n38477;
  assign n38479 = n8898 & n38478;
  assign n38480 = n8863 & n38479;
  assign n38481 = pi275 & ~n501;
  assign n38482 = n12872 & n38481;
  assign n38483 = n18049 & n38482;
  assign n38484 = n18053 & n38483;
  assign n38485 = n18047 & n38484;
  assign n38486 = n18080 & n38485;
  assign n38487 = ~n1172 & n38486;
  assign n38488 = ~n996 & n38487;
  assign n38489 = ~n2306 & n38488;
  assign n38490 = ~n500 & n38489;
  assign n38491 = n18038 & n38490;
  assign n38492 = n18037 & n38491;
  assign n38493 = n18088 & n38492;
  assign n38494 = n18106 & n38493;
  assign n38495 = n18035 & n38494;
  assign n38496 = n18134 & n38495;
  assign n38497 = ~n7236 & n38496;
  assign n38498 = ~n6137 & n38497;
  assign n38499 = n6193 & n38498;
  assign n38500 = n6134 & n38499;
  assign n38501 = ~n8867 & n38500;
  assign n38502 = ~n7235 & n38501;
  assign n38503 = n7296 & n38502;
  assign n38504 = n7231 & n38503;
  assign n38505 = ~n10027 & n38504;
  assign n38506 = ~n8866 & n38505;
  assign n38507 = n8898 & n38506;
  assign n38508 = n8863 & n38507;
  assign n38509 = ~n38480 & ~n38508;
  assign n38510 = ~n10788 & ~n38509;
  assign n38511 = ~n10026 & n38510;
  assign n38512 = n10072 & n38511;
  assign n38513 = n10021 & n38512;
  assign n38514 = ~n38452 & ~n38513;
  assign n38515 = ~n38449 & n38514;
  assign n38516 = ~n15278 & n35391;
  assign n38517 = ~n16216 & n38516;
  assign n38518 = n16939 & n38517;
  assign n38519 = ~n16937 & n38518;
  assign n38520 = n16944 & n38519;
  assign n38521 = n16936 & n38520;
  assign n38522 = ~n15167 & n35386;
  assign n38523 = ~n16216 & n38522;
  assign n38524 = ~n16220 & n38523;
  assign n38525 = ~n16466 & n38524;
  assign n38526 = n16476 & n38525;
  assign n38527 = ~n38521 & ~n38526;
  assign n38528 = n38515 & n38527;
  assign n38529 = ~n13764 & n35292;
  assign n38530 = ~n16216 & n38529;
  assign n38531 = ~n15465 & n38530;
  assign n38532 = ~n16209 & n38531;
  assign n38533 = n17086 & n38532;
  assign n38534 = n17133 & n38533;
  assign n38535 = n17122 & n38534;
  assign n38536 = ~n13726 & n35407;
  assign n38537 = ~n16216 & n38536;
  assign n38538 = ~n15419 & n38537;
  assign n38539 = n17086 & n38538;
  assign n38540 = n17094 & n38539;
  assign n38541 = n17083 & n38540;
  assign n38542 = ~n38535 & ~n38541;
  assign n38543 = n38528 & n38542;
  assign n38544 = n38445 & n38543;
  assign n38545 = n38411 & n38544;
  assign n38546 = pi259 & ~n16417;
  assign n38547 = ~n17766 & n38546;
  assign n38548 = ~n16216 & n38547;
  assign n38549 = ~n16215 & n38548;
  assign n38550 = n16222 & n38549;
  assign n38551 = n17637 & n38550;
  assign n38552 = n17629 & n38551;
  assign n38553 = n17765 & n38552;
  assign n38554 = n17874 & n38553;
  assign n38555 = pi171 & ~n8633;
  assign n38556 = ~n8455 & n38555;
  assign n38557 = ~n8834 & n38556;
  assign n38558 = ~n10002 & n38557;
  assign n38559 = ~n17152 & n38558;
  assign n38560 = ~n17151 & n38559;
  assign n38561 = ~n11297 & n38560;
  assign n38562 = ~n12240 & n38561;
  assign n38563 = ~n13135 & n38562;
  assign n38564 = ~n16216 & n38563;
  assign n38565 = ~n16215 & n38564;
  assign n38566 = n16222 & n38565;
  assign n38567 = n17163 & n38566;
  assign n38568 = n17167 & n38567;
  assign n38569 = n17150 & n38568;
  assign n38570 = n17192 & n38569;
  assign n38571 = ~n38554 & ~n38570;
  assign n38572 = ~n6401 & n27789;
  assign n38573 = ~n6784 & n38572;
  assign n38574 = ~n7158 & n38573;
  assign n38575 = ~n8250 & n38574;
  assign n38576 = ~n9414 & n38575;
  assign n38577 = ~n16957 & n38576;
  assign n38578 = ~n16956 & n38577;
  assign n38579 = ~n10667 & n38578;
  assign n38580 = ~n12083 & n38579;
  assign n38581 = ~n13644 & n38580;
  assign n38582 = ~n16216 & n38581;
  assign n38583 = ~n16215 & n38582;
  assign n38584 = n16222 & n38583;
  assign n38585 = n16971 & n38584;
  assign n38586 = n16975 & n38585;
  assign n38587 = n16955 & n38586;
  assign n38588 = n17000 & n38587;
  assign n38589 = ~n11042 & n35509;
  assign n38590 = ~n11188 & n38589;
  assign n38591 = ~n17378 & n38590;
  assign n38592 = ~n17377 & n38591;
  assign n38593 = ~n12380 & n38592;
  assign n38594 = ~n14045 & n38593;
  assign n38595 = ~n16216 & n38594;
  assign n38596 = ~n16215 & n38595;
  assign n38597 = n16222 & n38596;
  assign n38598 = n17387 & n38597;
  assign n38599 = n17391 & n38598;
  assign n38600 = n17376 & n38599;
  assign n38601 = n17416 & n38600;
  assign n38602 = ~n38588 & ~n38601;
  assign n38603 = n38571 & n38602;
  assign n38604 = ~n9763 & n35450;
  assign n38605 = ~n9929 & n38604;
  assign n38606 = ~n17263 & n38605;
  assign n38607 = ~n17262 & n38606;
  assign n38608 = ~n11266 & n38607;
  assign n38609 = ~n11588 & n38608;
  assign n38610 = ~n13859 & n38609;
  assign n38611 = ~n16216 & n38610;
  assign n38612 = ~n16215 & n38611;
  assign n38613 = n16222 & n38612;
  assign n38614 = n17273 & n38613;
  assign n38615 = n17277 & n38614;
  assign n38616 = n17261 & n38615;
  assign n38617 = n17302 & n38616;
  assign n38618 = pi123 & ~n5686;
  assign n38619 = ~n5349 & n38618;
  assign n38620 = ~n5808 & n38619;
  assign n38621 = ~n6056 & n38620;
  assign n38622 = ~n7073 & n38621;
  assign n38623 = ~n8179 & n38622;
  assign n38624 = ~n9344 & n38623;
  assign n38625 = ~n16418 & n38624;
  assign n38626 = ~n16361 & n38625;
  assign n38627 = ~n10594 & n38626;
  assign n38628 = ~n12005 & n38627;
  assign n38629 = ~n13558 & n38628;
  assign n38630 = ~n16216 & n38629;
  assign n38631 = ~n16215 & n38630;
  assign n38632 = n16432 & n38631;
  assign n38633 = n16435 & n38632;
  assign n38634 = n16439 & n38633;
  assign n38635 = n16305 & n38634;
  assign n38636 = n16464 & n38635;
  assign n38637 = ~n38617 & ~n38636;
  assign n38638 = ~n4460 & n35480;
  assign n38639 = ~n4817 & n38638;
  assign n38640 = ~n4902 & n38639;
  assign n38641 = ~n6001 & n38640;
  assign n38642 = ~n7014 & n38641;
  assign n38643 = ~n8114 & n38642;
  assign n38644 = ~n9276 & n38643;
  assign n38645 = ~n16486 & n38644;
  assign n38646 = ~n16485 & n38645;
  assign n38647 = ~n10523 & n38646;
  assign n38648 = ~n11928 & n38647;
  assign n38649 = ~n13479 & n38648;
  assign n38650 = ~n16216 & n38649;
  assign n38651 = ~n16220 & n38650;
  assign n38652 = n16503 & n38651;
  assign n38653 = n16506 & n38652;
  assign n38654 = n16510 & n38653;
  assign n38655 = n16484 & n38654;
  assign n38656 = n16535 & n38655;
  assign n38657 = pi059 & ~n1526;
  assign n38658 = ~n1556 & n38657;
  assign n38659 = ~n2242 & n38658;
  assign n38660 = ~n3095 & n38659;
  assign n38661 = ~n3997 & n38660;
  assign n38662 = ~n4003 & n38661;
  assign n38663 = ~n4837 & n38662;
  assign n38664 = ~n5822 & n38663;
  assign n38665 = ~n6820 & n38664;
  assign n38666 = ~n7785 & n38665;
  assign n38667 = ~n9027 & n38666;
  assign n38668 = ~n10245 & n38667;
  assign n38669 = ~n16748 & n38668;
  assign n38670 = ~n16747 & n38669;
  assign n38671 = ~n11536 & n38670;
  assign n38672 = ~n13036 & n38671;
  assign n38673 = ~n14653 & n38672;
  assign n38674 = ~n16746 & n38673;
  assign n38675 = ~n16745 & n38674;
  assign n38676 = n16770 & n38675;
  assign n38677 = n16773 & n38676;
  assign n38678 = n16777 & n38677;
  assign n38679 = n16744 & n38678;
  assign n38680 = n16802 & n38679;
  assign n38681 = ~n38656 & ~n38680;
  assign n38682 = n38637 & n38681;
  assign n38683 = ~n7505 & n23945;
  assign n38684 = ~n7869 & n38683;
  assign n38685 = ~n8346 & n38684;
  assign n38686 = ~n9485 & n38685;
  assign n38687 = ~n17018 & n38686;
  assign n38688 = ~n17017 & n38687;
  assign n38689 = ~n10741 & n38688;
  assign n38690 = ~n12158 & n38689;
  assign n38691 = ~n13693 & n38690;
  assign n38692 = ~n16216 & n38691;
  assign n38693 = ~n16215 & n38692;
  assign n38694 = n16222 & n38693;
  assign n38695 = n17031 & n38694;
  assign n38696 = n17035 & n38695;
  assign n38697 = n17016 & n38696;
  assign n38698 = n17060 & n38697;
  assign n38699 = ~n16216 & n35500;
  assign n38700 = ~n16215 & n38699;
  assign n38701 = n16222 & n38700;
  assign n38702 = n16225 & n38701;
  assign n38703 = n16229 & n38702;
  assign n38704 = n16214 & n38703;
  assign n38705 = n16297 & n38704;
  assign n38706 = ~n38698 & ~n38705;
  assign n38707 = pi075 & ~n2602;
  assign n38708 = ~n2783 & n38707;
  assign n38709 = ~n3066 & n38708;
  assign n38710 = ~n3983 & n38709;
  assign n38711 = ~n4003 & n38710;
  assign n38712 = ~n4024 & n38711;
  assign n38713 = ~n4999 & n38712;
  assign n38714 = ~n5827 & n38713;
  assign n38715 = ~n6893 & n38714;
  assign n38716 = ~n7890 & n38715;
  assign n38717 = ~n9131 & n38716;
  assign n38718 = ~n16617 & n38717;
  assign n38719 = ~n16616 & n38718;
  assign n38720 = ~n10278 & n38719;
  assign n38721 = ~n11662 & n38720;
  assign n38722 = ~n13191 & n38721;
  assign n38723 = ~n16615 & n38722;
  assign n38724 = ~n16614 & n38723;
  assign n38725 = n16636 & n38724;
  assign n38726 = n16639 & n38725;
  assign n38727 = n16643 & n38726;
  assign n38728 = n16613 & n38727;
  assign n38729 = n16668 & n38728;
  assign n38730 = pi235 & ~n14350;
  assign n38731 = ~n14381 & n38730;
  assign n38732 = ~n14519 & n38731;
  assign n38733 = ~n17537 & n38732;
  assign n38734 = ~n17536 & n38733;
  assign n38735 = ~n16216 & n38734;
  assign n38736 = ~n16215 & n38735;
  assign n38737 = n16222 & n38736;
  assign n38738 = n17544 & n38737;
  assign n38739 = n17547 & n38738;
  assign n38740 = n16214 & n38739;
  assign n38741 = n17572 & n38740;
  assign n38742 = ~n38729 & ~n38741;
  assign n38743 = n38706 & n38742;
  assign n38744 = n38682 & n38743;
  assign n38745 = n38603 & n38744;
  assign po140 = ~n38545 | ~n38745;
  assign n38747 = ~n3650 & n28036;
  assign n38748 = ~n3940 & n38747;
  assign n38749 = ~n4001 & n38748;
  assign n38750 = ~n5043 & n38749;
  assign n38751 = ~n5943 & n38750;
  assign n38752 = ~n6951 & n38751;
  assign n38753 = ~n8037 & n38752;
  assign n38754 = ~n9200 & n38753;
  assign n38755 = ~n16555 & n38754;
  assign n38756 = ~n16554 & n38755;
  assign n38757 = ~n10445 & n38756;
  assign n38758 = ~n11846 & n38757;
  assign n38759 = ~n13393 & n38758;
  assign n38760 = ~n16216 & n38759;
  assign n38761 = ~n16553 & n38760;
  assign n38762 = n16573 & n38761;
  assign n38763 = n16576 & n38762;
  assign n38764 = n16580 & n38763;
  assign n38765 = n16552 & n38764;
  assign n38766 = n16605 & n38765;
  assign n38767 = pi252 & ~n16144;
  assign n38768 = ~n16175 & n38767;
  assign n38769 = ~n16360 & n38768;
  assign n38770 = ~n17630 & n38769;
  assign n38771 = ~n16216 & n38770;
  assign n38772 = ~n16215 & n38771;
  assign n38773 = n16222 & n38772;
  assign n38774 = n17637 & n38773;
  assign n38775 = n17629 & n38774;
  assign n38776 = n17628 & n38775;
  assign n38777 = n17736 & n38776;
  assign n38778 = ~n38766 & ~n38777;
  assign n38779 = ~n780 & n27997;
  assign n38780 = ~n1372 & n38779;
  assign n38781 = ~n2243 & n38780;
  assign n38782 = ~n3104 & n38781;
  assign n38783 = ~n3971 & n38782;
  assign n38784 = ~n16682 & n38783;
  assign n38785 = ~n4872 & n38784;
  assign n38786 = ~n5801 & n38785;
  assign n38787 = ~n6739 & n38786;
  assign n38788 = ~n7807 & n38787;
  assign n38789 = ~n8989 & n38788;
  assign n38790 = ~n10273 & n38789;
  assign n38791 = ~n16680 & n38790;
  assign n38792 = ~n16679 & n38791;
  assign n38793 = ~n11499 & n38792;
  assign n38794 = ~n13076 & n38793;
  assign n38795 = ~n14698 & n38794;
  assign n38796 = ~n16678 & n38795;
  assign n38797 = ~n16677 & n38796;
  assign n38798 = n16704 & n38797;
  assign n38799 = n16707 & n38798;
  assign n38800 = n16711 & n38799;
  assign n38801 = n16676 & n38800;
  assign n38802 = n16736 & n38801;
  assign n38803 = pi220 & ~n12743;
  assign n38804 = ~n12773 & n38803;
  assign n38805 = ~n12902 & n38804;
  assign n38806 = ~n17419 & n38805;
  assign n38807 = ~n17418 & n38806;
  assign n38808 = ~n14009 & n38807;
  assign n38809 = ~n16216 & n38808;
  assign n38810 = ~n16215 & n38809;
  assign n38811 = n16222 & n38810;
  assign n38812 = n17427 & n38811;
  assign n38813 = n17431 & n38812;
  assign n38814 = n16214 & n38813;
  assign n38815 = n17456 & n38814;
  assign n38816 = ~n38802 & ~n38815;
  assign n38817 = n38778 & n38816;
  assign n38818 = ~n13906 & n35659;
  assign n38819 = ~n16216 & n38818;
  assign n38820 = ~n15586 & n38819;
  assign n38821 = ~n16208 & n38820;
  assign n38822 = n17257 & n38821;
  assign n38823 = n17328 & n38822;
  assign n38824 = n17342 & n38823;
  assign n38825 = ~n13820 & n35772;
  assign n38826 = ~n16216 & n38825;
  assign n38827 = ~n14741 & n38826;
  assign n38828 = ~n16209 & n38827;
  assign n38829 = ~n16211 & n38828;
  assign n38830 = n17238 & n38829;
  assign n38831 = n17232 & n38830;
  assign n38832 = n17225 & n38831;
  assign n38833 = ~n38824 & ~n38832;
  assign n38834 = ~n14073 & n35764;
  assign n38835 = ~n16216 & n38834;
  assign n38836 = ~n15616 & n38835;
  assign n38837 = ~n16224 & n38836;
  assign n38838 = n17086 & n38837;
  assign n38839 = n17351 & n38838;
  assign n38840 = n17350 & n38839;
  assign n38841 = n17370 & n38840;
  assign n38842 = ~n13093 & n32925;
  assign n38843 = ~n16216 & n38842;
  assign n38844 = ~n16215 & n38843;
  assign n38845 = n16222 & n38844;
  assign n38846 = n17516 & n38845;
  assign n38847 = n16214 & n38846;
  assign n38848 = n17512 & n38847;
  assign n38849 = n17534 & n38848;
  assign n38850 = ~n38841 & ~n38849;
  assign n38851 = n38833 & n38850;
  assign n38852 = ~n15075 & n35681;
  assign n38853 = ~n16216 & n38852;
  assign n38854 = ~n16537 & n38853;
  assign n38855 = n16544 & n38854;
  assign n38856 = ~n16831 & n35685;
  assign n38857 = ~n16829 & n38856;
  assign n38858 = n16836 & n38857;
  assign n38859 = pi268 & ~n501;
  assign n38860 = n12872 & n38859;
  assign n38861 = n17949 & n38860;
  assign n38862 = n17954 & n38861;
  assign n38863 = n17947 & n38862;
  assign n38864 = n17982 & n38863;
  assign n38865 = ~n1172 & n38864;
  assign n38866 = ~n996 & n38865;
  assign n38867 = ~n2306 & n38866;
  assign n38868 = ~n500 & n38867;
  assign n38869 = n17940 & n38868;
  assign n38870 = n17991 & n38869;
  assign n38871 = n17938 & n38870;
  assign n38872 = n17929 & n38871;
  assign n38873 = n17921 & n38872;
  assign n38874 = n18029 & n38873;
  assign n38875 = ~n7236 & n38874;
  assign n38876 = ~n6137 & n38875;
  assign n38877 = n6193 & n38876;
  assign n38878 = n6134 & n38877;
  assign n38879 = ~n8867 & n38878;
  assign n38880 = ~n7235 & n38879;
  assign n38881 = n7296 & n38880;
  assign n38882 = n7231 & n38881;
  assign n38883 = ~n10027 & n38882;
  assign n38884 = ~n8866 & n38883;
  assign n38885 = n8898 & n38884;
  assign n38886 = n8863 & n38885;
  assign n38887 = pi276 & ~n501;
  assign n38888 = n12872 & n38887;
  assign n38889 = n18049 & n38888;
  assign n38890 = n18053 & n38889;
  assign n38891 = n18047 & n38890;
  assign n38892 = n18080 & n38891;
  assign n38893 = ~n1172 & n38892;
  assign n38894 = ~n996 & n38893;
  assign n38895 = ~n2306 & n38894;
  assign n38896 = ~n500 & n38895;
  assign n38897 = n18038 & n38896;
  assign n38898 = n18037 & n38897;
  assign n38899 = n18088 & n38898;
  assign n38900 = n18106 & n38899;
  assign n38901 = n18035 & n38900;
  assign n38902 = n18134 & n38901;
  assign n38903 = ~n7236 & n38902;
  assign n38904 = ~n6137 & n38903;
  assign n38905 = n6193 & n38904;
  assign n38906 = n6134 & n38905;
  assign n38907 = ~n8867 & n38906;
  assign n38908 = ~n7235 & n38907;
  assign n38909 = n7296 & n38908;
  assign n38910 = n7231 & n38909;
  assign n38911 = ~n10027 & n38910;
  assign n38912 = ~n8866 & n38911;
  assign n38913 = n8898 & n38912;
  assign n38914 = n8863 & n38913;
  assign n38915 = ~n38886 & ~n38914;
  assign n38916 = ~n10788 & ~n38915;
  assign n38917 = ~n10026 & n38916;
  assign n38918 = n10072 & n38917;
  assign n38919 = n10021 & n38918;
  assign n38920 = ~n38858 & ~n38919;
  assign n38921 = ~n38855 & n38920;
  assign n38922 = ~n15278 & n35756;
  assign n38923 = ~n16216 & n38922;
  assign n38924 = n16939 & n38923;
  assign n38925 = ~n16937 & n38924;
  assign n38926 = n16944 & n38925;
  assign n38927 = n16936 & n38926;
  assign n38928 = ~n15167 & n35751;
  assign n38929 = ~n16216 & n38928;
  assign n38930 = ~n16220 & n38929;
  assign n38931 = ~n16466 & n38930;
  assign n38932 = n16476 & n38931;
  assign n38933 = ~n38927 & ~n38932;
  assign n38934 = n38921 & n38933;
  assign n38935 = ~n13764 & n35666;
  assign n38936 = ~n16216 & n38935;
  assign n38937 = ~n15465 & n38936;
  assign n38938 = ~n16209 & n38937;
  assign n38939 = n17086 & n38938;
  assign n38940 = n17133 & n38939;
  assign n38941 = n17122 & n38940;
  assign n38942 = ~n13726 & n35673;
  assign n38943 = ~n16216 & n38942;
  assign n38944 = ~n15419 & n38943;
  assign n38945 = n17086 & n38944;
  assign n38946 = n17094 & n38945;
  assign n38947 = n17083 & n38946;
  assign n38948 = ~n38941 & ~n38947;
  assign n38949 = n38934 & n38948;
  assign n38950 = n38851 & n38949;
  assign n38951 = n38817 & n38950;
  assign n38952 = pi260 & ~n16417;
  assign n38953 = ~n17766 & n38952;
  assign n38954 = ~n16216 & n38953;
  assign n38955 = ~n16215 & n38954;
  assign n38956 = n16222 & n38955;
  assign n38957 = n17637 & n38956;
  assign n38958 = n17629 & n38957;
  assign n38959 = n17765 & n38958;
  assign n38960 = n17874 & n38959;
  assign n38961 = pi172 & ~n8633;
  assign n38962 = ~n8455 & n38961;
  assign n38963 = ~n8834 & n38962;
  assign n38964 = ~n10002 & n38963;
  assign n38965 = ~n17152 & n38964;
  assign n38966 = ~n17151 & n38965;
  assign n38967 = ~n11297 & n38966;
  assign n38968 = ~n12240 & n38967;
  assign n38969 = ~n13135 & n38968;
  assign n38970 = ~n16216 & n38969;
  assign n38971 = ~n16215 & n38970;
  assign n38972 = n16222 & n38971;
  assign n38973 = n17163 & n38972;
  assign n38974 = n17167 & n38973;
  assign n38975 = n17150 & n38974;
  assign n38976 = n17192 & n38975;
  assign n38977 = ~n38960 & ~n38976;
  assign n38978 = ~n6401 & n28055;
  assign n38979 = ~n6784 & n38978;
  assign n38980 = ~n7158 & n38979;
  assign n38981 = ~n8250 & n38980;
  assign n38982 = ~n9414 & n38981;
  assign n38983 = ~n16957 & n38982;
  assign n38984 = ~n16956 & n38983;
  assign n38985 = ~n10667 & n38984;
  assign n38986 = ~n12083 & n38985;
  assign n38987 = ~n13644 & n38986;
  assign n38988 = ~n16216 & n38987;
  assign n38989 = ~n16215 & n38988;
  assign n38990 = n16222 & n38989;
  assign n38991 = n16971 & n38990;
  assign n38992 = n16975 & n38991;
  assign n38993 = n16955 & n38992;
  assign n38994 = n17000 & n38993;
  assign n38995 = ~n11042 & n35632;
  assign n38996 = ~n11188 & n38995;
  assign n38997 = ~n17378 & n38996;
  assign n38998 = ~n17377 & n38997;
  assign n38999 = ~n12380 & n38998;
  assign n39000 = ~n14045 & n38999;
  assign n39001 = ~n16216 & n39000;
  assign n39002 = ~n16215 & n39001;
  assign n39003 = n16222 & n39002;
  assign n39004 = n17387 & n39003;
  assign n39005 = n17391 & n39004;
  assign n39006 = n17376 & n39005;
  assign n39007 = n17416 & n39006;
  assign n39008 = ~n38994 & ~n39007;
  assign n39009 = n38977 & n39008;
  assign n39010 = ~n9763 & n35822;
  assign n39011 = ~n9929 & n39010;
  assign n39012 = ~n17263 & n39011;
  assign n39013 = ~n17262 & n39012;
  assign n39014 = ~n11266 & n39013;
  assign n39015 = ~n11588 & n39014;
  assign n39016 = ~n13859 & n39015;
  assign n39017 = ~n16216 & n39016;
  assign n39018 = ~n16215 & n39017;
  assign n39019 = n16222 & n39018;
  assign n39020 = n17273 & n39019;
  assign n39021 = n17277 & n39020;
  assign n39022 = n17261 & n39021;
  assign n39023 = n17302 & n39022;
  assign n39024 = pi124 & ~n5686;
  assign n39025 = ~n5349 & n39024;
  assign n39026 = ~n5808 & n39025;
  assign n39027 = ~n6056 & n39026;
  assign n39028 = ~n7073 & n39027;
  assign n39029 = ~n8179 & n39028;
  assign n39030 = ~n9344 & n39029;
  assign n39031 = ~n16418 & n39030;
  assign n39032 = ~n16361 & n39031;
  assign n39033 = ~n10594 & n39032;
  assign n39034 = ~n12005 & n39033;
  assign n39035 = ~n13558 & n39034;
  assign n39036 = ~n16216 & n39035;
  assign n39037 = ~n16215 & n39036;
  assign n39038 = n16432 & n39037;
  assign n39039 = n16435 & n39038;
  assign n39040 = n16439 & n39039;
  assign n39041 = n16305 & n39040;
  assign n39042 = n16464 & n39041;
  assign n39043 = ~n39023 & ~n39042;
  assign n39044 = ~n4460 & n35838;
  assign n39045 = ~n4817 & n39044;
  assign n39046 = ~n4902 & n39045;
  assign n39047 = ~n6001 & n39046;
  assign n39048 = ~n7014 & n39047;
  assign n39049 = ~n8114 & n39048;
  assign n39050 = ~n9276 & n39049;
  assign n39051 = ~n16486 & n39050;
  assign n39052 = ~n16485 & n39051;
  assign n39053 = ~n10523 & n39052;
  assign n39054 = ~n11928 & n39053;
  assign n39055 = ~n13479 & n39054;
  assign n39056 = ~n16216 & n39055;
  assign n39057 = ~n16220 & n39056;
  assign n39058 = n16503 & n39057;
  assign n39059 = n16506 & n39058;
  assign n39060 = n16510 & n39059;
  assign n39061 = n16484 & n39060;
  assign n39062 = n16535 & n39061;
  assign n39063 = pi060 & ~n1526;
  assign n39064 = ~n1556 & n39063;
  assign n39065 = ~n2242 & n39064;
  assign n39066 = ~n3095 & n39065;
  assign n39067 = ~n3997 & n39066;
  assign n39068 = ~n4003 & n39067;
  assign n39069 = ~n4837 & n39068;
  assign n39070 = ~n5822 & n39069;
  assign n39071 = ~n6820 & n39070;
  assign n39072 = ~n7785 & n39071;
  assign n39073 = ~n9027 & n39072;
  assign n39074 = ~n10245 & n39073;
  assign n39075 = ~n16748 & n39074;
  assign n39076 = ~n16747 & n39075;
  assign n39077 = ~n11536 & n39076;
  assign n39078 = ~n13036 & n39077;
  assign n39079 = ~n14653 & n39078;
  assign n39080 = ~n16746 & n39079;
  assign n39081 = ~n16745 & n39080;
  assign n39082 = n16770 & n39081;
  assign n39083 = n16773 & n39082;
  assign n39084 = n16777 & n39083;
  assign n39085 = n16744 & n39084;
  assign n39086 = n16802 & n39085;
  assign n39087 = ~n39062 & ~n39086;
  assign n39088 = n39043 & n39087;
  assign n39089 = ~n7505 & n24206;
  assign n39090 = ~n7869 & n39089;
  assign n39091 = ~n8346 & n39090;
  assign n39092 = ~n9485 & n39091;
  assign n39093 = ~n17018 & n39092;
  assign n39094 = ~n17017 & n39093;
  assign n39095 = ~n10741 & n39094;
  assign n39096 = ~n12158 & n39095;
  assign n39097 = ~n13693 & n39096;
  assign n39098 = ~n16216 & n39097;
  assign n39099 = ~n16215 & n39098;
  assign n39100 = n16222 & n39099;
  assign n39101 = n17031 & n39100;
  assign n39102 = n17035 & n39101;
  assign n39103 = n17016 & n39102;
  assign n39104 = n17060 & n39103;
  assign n39105 = ~n16216 & n35622;
  assign n39106 = ~n16215 & n39105;
  assign n39107 = n16222 & n39106;
  assign n39108 = n16225 & n39107;
  assign n39109 = n16229 & n39108;
  assign n39110 = n16214 & n39109;
  assign n39111 = n16297 & n39110;
  assign n39112 = ~n39104 & ~n39111;
  assign n39113 = pi076 & ~n2602;
  assign n39114 = ~n2783 & n39113;
  assign n39115 = ~n3066 & n39114;
  assign n39116 = ~n3983 & n39115;
  assign n39117 = ~n4003 & n39116;
  assign n39118 = ~n4024 & n39117;
  assign n39119 = ~n4999 & n39118;
  assign n39120 = ~n5827 & n39119;
  assign n39121 = ~n6893 & n39120;
  assign n39122 = ~n7890 & n39121;
  assign n39123 = ~n9131 & n39122;
  assign n39124 = ~n16617 & n39123;
  assign n39125 = ~n16616 & n39124;
  assign n39126 = ~n10278 & n39125;
  assign n39127 = ~n11662 & n39126;
  assign n39128 = ~n13191 & n39127;
  assign n39129 = ~n16615 & n39128;
  assign n39130 = ~n16614 & n39129;
  assign n39131 = n16636 & n39130;
  assign n39132 = n16639 & n39131;
  assign n39133 = n16643 & n39132;
  assign n39134 = n16613 & n39133;
  assign n39135 = n16668 & n39134;
  assign n39136 = pi236 & ~n14350;
  assign n39137 = ~n14381 & n39136;
  assign n39138 = ~n14519 & n39137;
  assign n39139 = ~n17537 & n39138;
  assign n39140 = ~n17536 & n39139;
  assign n39141 = ~n16216 & n39140;
  assign n39142 = ~n16215 & n39141;
  assign n39143 = n16222 & n39142;
  assign n39144 = n17544 & n39143;
  assign n39145 = n17547 & n39144;
  assign n39146 = n16214 & n39145;
  assign n39147 = n17572 & n39146;
  assign n39148 = ~n39135 & ~n39147;
  assign n39149 = n39112 & n39148;
  assign n39150 = n39088 & n39149;
  assign n39151 = n39009 & n39150;
  assign po141 = ~n38951 | ~n39151;
  assign n39153 = ~n3650 & n28302;
  assign n39154 = ~n3940 & n39153;
  assign n39155 = ~n4001 & n39154;
  assign n39156 = ~n5043 & n39155;
  assign n39157 = ~n5943 & n39156;
  assign n39158 = ~n6951 & n39157;
  assign n39159 = ~n8037 & n39158;
  assign n39160 = ~n9200 & n39159;
  assign n39161 = ~n16555 & n39160;
  assign n39162 = ~n16554 & n39161;
  assign n39163 = ~n10445 & n39162;
  assign n39164 = ~n11846 & n39163;
  assign n39165 = ~n13393 & n39164;
  assign n39166 = ~n16216 & n39165;
  assign n39167 = ~n16553 & n39166;
  assign n39168 = n16573 & n39167;
  assign n39169 = n16576 & n39168;
  assign n39170 = n16580 & n39169;
  assign n39171 = n16552 & n39170;
  assign n39172 = n16605 & n39171;
  assign n39173 = pi253 & ~n16144;
  assign n39174 = ~n16175 & n39173;
  assign n39175 = ~n16360 & n39174;
  assign n39176 = ~n17630 & n39175;
  assign n39177 = ~n16216 & n39176;
  assign n39178 = ~n16215 & n39177;
  assign n39179 = n16222 & n39178;
  assign n39180 = n17637 & n39179;
  assign n39181 = n17629 & n39180;
  assign n39182 = n17628 & n39181;
  assign n39183 = n17736 & n39182;
  assign n39184 = ~n39172 & ~n39183;
  assign n39185 = ~n780 & n28263;
  assign n39186 = ~n1372 & n39185;
  assign n39187 = ~n2243 & n39186;
  assign n39188 = ~n3104 & n39187;
  assign n39189 = ~n3971 & n39188;
  assign n39190 = ~n16682 & n39189;
  assign n39191 = ~n4872 & n39190;
  assign n39192 = ~n5801 & n39191;
  assign n39193 = ~n6739 & n39192;
  assign n39194 = ~n7807 & n39193;
  assign n39195 = ~n8989 & n39194;
  assign n39196 = ~n10273 & n39195;
  assign n39197 = ~n16680 & n39196;
  assign n39198 = ~n16679 & n39197;
  assign n39199 = ~n11499 & n39198;
  assign n39200 = ~n13076 & n39199;
  assign n39201 = ~n14698 & n39200;
  assign n39202 = ~n16678 & n39201;
  assign n39203 = ~n16677 & n39202;
  assign n39204 = n16704 & n39203;
  assign n39205 = n16707 & n39204;
  assign n39206 = n16711 & n39205;
  assign n39207 = n16676 & n39206;
  assign n39208 = n16736 & n39207;
  assign n39209 = pi221 & ~n12743;
  assign n39210 = ~n12773 & n39209;
  assign n39211 = ~n12902 & n39210;
  assign n39212 = ~n17419 & n39211;
  assign n39213 = ~n17418 & n39212;
  assign n39214 = ~n14009 & n39213;
  assign n39215 = ~n16216 & n39214;
  assign n39216 = ~n16215 & n39215;
  assign n39217 = n16222 & n39216;
  assign n39218 = n17427 & n39217;
  assign n39219 = n17431 & n39218;
  assign n39220 = n16214 & n39219;
  assign n39221 = n17456 & n39220;
  assign n39222 = ~n39208 & ~n39221;
  assign n39223 = n39184 & n39222;
  assign n39224 = ~n13906 & n36031;
  assign n39225 = ~n16216 & n39224;
  assign n39226 = ~n15586 & n39225;
  assign n39227 = ~n16208 & n39226;
  assign n39228 = n17257 & n39227;
  assign n39229 = n17328 & n39228;
  assign n39230 = n17342 & n39229;
  assign n39231 = ~n13820 & n36144;
  assign n39232 = ~n16216 & n39231;
  assign n39233 = ~n14741 & n39232;
  assign n39234 = ~n16209 & n39233;
  assign n39235 = ~n16211 & n39234;
  assign n39236 = n17238 & n39235;
  assign n39237 = n17232 & n39236;
  assign n39238 = n17225 & n39237;
  assign n39239 = ~n39230 & ~n39238;
  assign n39240 = ~n14073 & n36136;
  assign n39241 = ~n16216 & n39240;
  assign n39242 = ~n15616 & n39241;
  assign n39243 = ~n16224 & n39242;
  assign n39244 = n17086 & n39243;
  assign n39245 = n17351 & n39244;
  assign n39246 = n17350 & n39245;
  assign n39247 = n17370 & n39246;
  assign n39248 = ~n13093 & n33250;
  assign n39249 = ~n16216 & n39248;
  assign n39250 = ~n16215 & n39249;
  assign n39251 = n16222 & n39250;
  assign n39252 = n17516 & n39251;
  assign n39253 = n16214 & n39252;
  assign n39254 = n17512 & n39253;
  assign n39255 = n17534 & n39254;
  assign n39256 = ~n39247 & ~n39255;
  assign n39257 = n39239 & n39256;
  assign n39258 = ~n15075 & n36053;
  assign n39259 = ~n16216 & n39258;
  assign n39260 = ~n16537 & n39259;
  assign n39261 = n16544 & n39260;
  assign n39262 = ~n16831 & n36057;
  assign n39263 = ~n16829 & n39262;
  assign n39264 = n16836 & n39263;
  assign n39265 = pi269 & ~n501;
  assign n39266 = n12872 & n39265;
  assign n39267 = n17949 & n39266;
  assign n39268 = n17954 & n39267;
  assign n39269 = n17947 & n39268;
  assign n39270 = n17982 & n39269;
  assign n39271 = ~n1172 & n39270;
  assign n39272 = ~n996 & n39271;
  assign n39273 = ~n2306 & n39272;
  assign n39274 = ~n500 & n39273;
  assign n39275 = n17940 & n39274;
  assign n39276 = n17991 & n39275;
  assign n39277 = n17938 & n39276;
  assign n39278 = n17929 & n39277;
  assign n39279 = n17921 & n39278;
  assign n39280 = n18029 & n39279;
  assign n39281 = ~n7236 & n39280;
  assign n39282 = ~n6137 & n39281;
  assign n39283 = n6193 & n39282;
  assign n39284 = n6134 & n39283;
  assign n39285 = ~n8867 & n39284;
  assign n39286 = ~n7235 & n39285;
  assign n39287 = n7296 & n39286;
  assign n39288 = n7231 & n39287;
  assign n39289 = ~n10027 & n39288;
  assign n39290 = ~n8866 & n39289;
  assign n39291 = n8898 & n39290;
  assign n39292 = n8863 & n39291;
  assign n39293 = pi277 & ~n501;
  assign n39294 = n12872 & n39293;
  assign n39295 = n18049 & n39294;
  assign n39296 = n18053 & n39295;
  assign n39297 = n18047 & n39296;
  assign n39298 = n18080 & n39297;
  assign n39299 = ~n1172 & n39298;
  assign n39300 = ~n996 & n39299;
  assign n39301 = ~n2306 & n39300;
  assign n39302 = ~n500 & n39301;
  assign n39303 = n18038 & n39302;
  assign n39304 = n18037 & n39303;
  assign n39305 = n18088 & n39304;
  assign n39306 = n18106 & n39305;
  assign n39307 = n18035 & n39306;
  assign n39308 = n18134 & n39307;
  assign n39309 = ~n7236 & n39308;
  assign n39310 = ~n6137 & n39309;
  assign n39311 = n6193 & n39310;
  assign n39312 = n6134 & n39311;
  assign n39313 = ~n8867 & n39312;
  assign n39314 = ~n7235 & n39313;
  assign n39315 = n7296 & n39314;
  assign n39316 = n7231 & n39315;
  assign n39317 = ~n10027 & n39316;
  assign n39318 = ~n8866 & n39317;
  assign n39319 = n8898 & n39318;
  assign n39320 = n8863 & n39319;
  assign n39321 = ~n39292 & ~n39320;
  assign n39322 = ~n10788 & ~n39321;
  assign n39323 = ~n10026 & n39322;
  assign n39324 = n10072 & n39323;
  assign n39325 = n10021 & n39324;
  assign n39326 = ~n39264 & ~n39325;
  assign n39327 = ~n39261 & n39326;
  assign n39328 = ~n15278 & n36128;
  assign n39329 = ~n16216 & n39328;
  assign n39330 = n16939 & n39329;
  assign n39331 = ~n16937 & n39330;
  assign n39332 = n16944 & n39331;
  assign n39333 = n16936 & n39332;
  assign n39334 = ~n15167 & n36123;
  assign n39335 = ~n16216 & n39334;
  assign n39336 = ~n16220 & n39335;
  assign n39337 = ~n16466 & n39336;
  assign n39338 = n16476 & n39337;
  assign n39339 = ~n39333 & ~n39338;
  assign n39340 = n39327 & n39339;
  assign n39341 = ~n13764 & n36038;
  assign n39342 = ~n16216 & n39341;
  assign n39343 = ~n15465 & n39342;
  assign n39344 = ~n16209 & n39343;
  assign n39345 = n17086 & n39344;
  assign n39346 = n17133 & n39345;
  assign n39347 = n17122 & n39346;
  assign n39348 = ~n13726 & n36045;
  assign n39349 = ~n16216 & n39348;
  assign n39350 = ~n15419 & n39349;
  assign n39351 = n17086 & n39350;
  assign n39352 = n17094 & n39351;
  assign n39353 = n17083 & n39352;
  assign n39354 = ~n39347 & ~n39353;
  assign n39355 = n39340 & n39354;
  assign n39356 = n39257 & n39355;
  assign n39357 = n39223 & n39356;
  assign n39358 = pi261 & ~n16417;
  assign n39359 = ~n17766 & n39358;
  assign n39360 = ~n16216 & n39359;
  assign n39361 = ~n16215 & n39360;
  assign n39362 = n16222 & n39361;
  assign n39363 = n17637 & n39362;
  assign n39364 = n17629 & n39363;
  assign n39365 = n17765 & n39364;
  assign n39366 = n17874 & n39365;
  assign n39367 = pi173 & ~n8633;
  assign n39368 = ~n8455 & n39367;
  assign n39369 = ~n8834 & n39368;
  assign n39370 = ~n10002 & n39369;
  assign n39371 = ~n17152 & n39370;
  assign n39372 = ~n17151 & n39371;
  assign n39373 = ~n11297 & n39372;
  assign n39374 = ~n12240 & n39373;
  assign n39375 = ~n13135 & n39374;
  assign n39376 = ~n16216 & n39375;
  assign n39377 = ~n16215 & n39376;
  assign n39378 = n16222 & n39377;
  assign n39379 = n17163 & n39378;
  assign n39380 = n17167 & n39379;
  assign n39381 = n17150 & n39380;
  assign n39382 = n17192 & n39381;
  assign n39383 = ~n39366 & ~n39382;
  assign n39384 = ~n6401 & n28321;
  assign n39385 = ~n6784 & n39384;
  assign n39386 = ~n7158 & n39385;
  assign n39387 = ~n8250 & n39386;
  assign n39388 = ~n9414 & n39387;
  assign n39389 = ~n16957 & n39388;
  assign n39390 = ~n16956 & n39389;
  assign n39391 = ~n10667 & n39390;
  assign n39392 = ~n12083 & n39391;
  assign n39393 = ~n13644 & n39392;
  assign n39394 = ~n16216 & n39393;
  assign n39395 = ~n16215 & n39394;
  assign n39396 = n16222 & n39395;
  assign n39397 = n16971 & n39396;
  assign n39398 = n16975 & n39397;
  assign n39399 = n16955 & n39398;
  assign n39400 = n17000 & n39399;
  assign n39401 = ~n11042 & n36004;
  assign n39402 = ~n11188 & n39401;
  assign n39403 = ~n17378 & n39402;
  assign n39404 = ~n17377 & n39403;
  assign n39405 = ~n12380 & n39404;
  assign n39406 = ~n14045 & n39405;
  assign n39407 = ~n16216 & n39406;
  assign n39408 = ~n16215 & n39407;
  assign n39409 = n16222 & n39408;
  assign n39410 = n17387 & n39409;
  assign n39411 = n17391 & n39410;
  assign n39412 = n17376 & n39411;
  assign n39413 = n17416 & n39412;
  assign n39414 = ~n39400 & ~n39413;
  assign n39415 = n39383 & n39414;
  assign n39416 = ~n9763 & n36194;
  assign n39417 = ~n9929 & n39416;
  assign n39418 = ~n17263 & n39417;
  assign n39419 = ~n17262 & n39418;
  assign n39420 = ~n11266 & n39419;
  assign n39421 = ~n11588 & n39420;
  assign n39422 = ~n13859 & n39421;
  assign n39423 = ~n16216 & n39422;
  assign n39424 = ~n16215 & n39423;
  assign n39425 = n16222 & n39424;
  assign n39426 = n17273 & n39425;
  assign n39427 = n17277 & n39426;
  assign n39428 = n17261 & n39427;
  assign n39429 = n17302 & n39428;
  assign n39430 = pi125 & ~n5686;
  assign n39431 = ~n5349 & n39430;
  assign n39432 = ~n5808 & n39431;
  assign n39433 = ~n6056 & n39432;
  assign n39434 = ~n7073 & n39433;
  assign n39435 = ~n8179 & n39434;
  assign n39436 = ~n9344 & n39435;
  assign n39437 = ~n16418 & n39436;
  assign n39438 = ~n16361 & n39437;
  assign n39439 = ~n10594 & n39438;
  assign n39440 = ~n12005 & n39439;
  assign n39441 = ~n13558 & n39440;
  assign n39442 = ~n16216 & n39441;
  assign n39443 = ~n16215 & n39442;
  assign n39444 = n16432 & n39443;
  assign n39445 = n16435 & n39444;
  assign n39446 = n16439 & n39445;
  assign n39447 = n16305 & n39446;
  assign n39448 = n16464 & n39447;
  assign n39449 = ~n39429 & ~n39448;
  assign n39450 = ~n4460 & n36210;
  assign n39451 = ~n4817 & n39450;
  assign n39452 = ~n4902 & n39451;
  assign n39453 = ~n6001 & n39452;
  assign n39454 = ~n7014 & n39453;
  assign n39455 = ~n8114 & n39454;
  assign n39456 = ~n9276 & n39455;
  assign n39457 = ~n16486 & n39456;
  assign n39458 = ~n16485 & n39457;
  assign n39459 = ~n10523 & n39458;
  assign n39460 = ~n11928 & n39459;
  assign n39461 = ~n13479 & n39460;
  assign n39462 = ~n16216 & n39461;
  assign n39463 = ~n16220 & n39462;
  assign n39464 = n16503 & n39463;
  assign n39465 = n16506 & n39464;
  assign n39466 = n16510 & n39465;
  assign n39467 = n16484 & n39466;
  assign n39468 = n16535 & n39467;
  assign n39469 = pi061 & ~n1526;
  assign n39470 = ~n1556 & n39469;
  assign n39471 = ~n2242 & n39470;
  assign n39472 = ~n3095 & n39471;
  assign n39473 = ~n3997 & n39472;
  assign n39474 = ~n4003 & n39473;
  assign n39475 = ~n4837 & n39474;
  assign n39476 = ~n5822 & n39475;
  assign n39477 = ~n6820 & n39476;
  assign n39478 = ~n7785 & n39477;
  assign n39479 = ~n9027 & n39478;
  assign n39480 = ~n10245 & n39479;
  assign n39481 = ~n16748 & n39480;
  assign n39482 = ~n16747 & n39481;
  assign n39483 = ~n11536 & n39482;
  assign n39484 = ~n13036 & n39483;
  assign n39485 = ~n14653 & n39484;
  assign n39486 = ~n16746 & n39485;
  assign n39487 = ~n16745 & n39486;
  assign n39488 = n16770 & n39487;
  assign n39489 = n16773 & n39488;
  assign n39490 = n16777 & n39489;
  assign n39491 = n16744 & n39490;
  assign n39492 = n16802 & n39491;
  assign n39493 = ~n39468 & ~n39492;
  assign n39494 = n39449 & n39493;
  assign n39495 = ~n7505 & n24399;
  assign n39496 = ~n7869 & n39495;
  assign n39497 = ~n8346 & n39496;
  assign n39498 = ~n9485 & n39497;
  assign n39499 = ~n17018 & n39498;
  assign n39500 = ~n17017 & n39499;
  assign n39501 = ~n10741 & n39500;
  assign n39502 = ~n12158 & n39501;
  assign n39503 = ~n13693 & n39502;
  assign n39504 = ~n16216 & n39503;
  assign n39505 = ~n16215 & n39504;
  assign n39506 = n16222 & n39505;
  assign n39507 = n17031 & n39506;
  assign n39508 = n17035 & n39507;
  assign n39509 = n17016 & n39508;
  assign n39510 = n17060 & n39509;
  assign n39511 = ~n16216 & n35994;
  assign n39512 = ~n16215 & n39511;
  assign n39513 = n16222 & n39512;
  assign n39514 = n16225 & n39513;
  assign n39515 = n16229 & n39514;
  assign n39516 = n16214 & n39515;
  assign n39517 = n16297 & n39516;
  assign n39518 = ~n39510 & ~n39517;
  assign n39519 = pi077 & ~n2602;
  assign n39520 = ~n2783 & n39519;
  assign n39521 = ~n3066 & n39520;
  assign n39522 = ~n3983 & n39521;
  assign n39523 = ~n4003 & n39522;
  assign n39524 = ~n4024 & n39523;
  assign n39525 = ~n4999 & n39524;
  assign n39526 = ~n5827 & n39525;
  assign n39527 = ~n6893 & n39526;
  assign n39528 = ~n7890 & n39527;
  assign n39529 = ~n9131 & n39528;
  assign n39530 = ~n16617 & n39529;
  assign n39531 = ~n16616 & n39530;
  assign n39532 = ~n10278 & n39531;
  assign n39533 = ~n11662 & n39532;
  assign n39534 = ~n13191 & n39533;
  assign n39535 = ~n16615 & n39534;
  assign n39536 = ~n16614 & n39535;
  assign n39537 = n16636 & n39536;
  assign n39538 = n16639 & n39537;
  assign n39539 = n16643 & n39538;
  assign n39540 = n16613 & n39539;
  assign n39541 = n16668 & n39540;
  assign n39542 = pi237 & ~n14350;
  assign n39543 = ~n14381 & n39542;
  assign n39544 = ~n14519 & n39543;
  assign n39545 = ~n17537 & n39544;
  assign n39546 = ~n17536 & n39545;
  assign n39547 = ~n16216 & n39546;
  assign n39548 = ~n16215 & n39547;
  assign n39549 = n16222 & n39548;
  assign n39550 = n17544 & n39549;
  assign n39551 = n17547 & n39550;
  assign n39552 = n16214 & n39551;
  assign n39553 = n17572 & n39552;
  assign n39554 = ~n39541 & ~n39553;
  assign n39555 = n39518 & n39554;
  assign n39556 = n39494 & n39555;
  assign n39557 = n39415 & n39556;
  assign po142 = ~n39357 | ~n39557;
  assign n39559 = ~n3650 & n28568;
  assign n39560 = ~n3940 & n39559;
  assign n39561 = ~n4001 & n39560;
  assign n39562 = ~n5043 & n39561;
  assign n39563 = ~n5943 & n39562;
  assign n39564 = ~n6951 & n39563;
  assign n39565 = ~n8037 & n39564;
  assign n39566 = ~n9200 & n39565;
  assign n39567 = ~n16555 & n39566;
  assign n39568 = ~n16554 & n39567;
  assign n39569 = ~n10445 & n39568;
  assign n39570 = ~n11846 & n39569;
  assign n39571 = ~n13393 & n39570;
  assign n39572 = ~n16216 & n39571;
  assign n39573 = ~n16553 & n39572;
  assign n39574 = n16573 & n39573;
  assign n39575 = n16576 & n39574;
  assign n39576 = n16580 & n39575;
  assign n39577 = n16552 & n39576;
  assign n39578 = n16605 & n39577;
  assign n39579 = pi254 & ~n16144;
  assign n39580 = ~n16175 & n39579;
  assign n39581 = ~n16360 & n39580;
  assign n39582 = ~n17630 & n39581;
  assign n39583 = ~n16216 & n39582;
  assign n39584 = ~n16215 & n39583;
  assign n39585 = n16222 & n39584;
  assign n39586 = n17637 & n39585;
  assign n39587 = n17629 & n39586;
  assign n39588 = n17628 & n39587;
  assign n39589 = n17736 & n39588;
  assign n39590 = ~n39578 & ~n39589;
  assign n39591 = ~n780 & n28529;
  assign n39592 = ~n1372 & n39591;
  assign n39593 = ~n2243 & n39592;
  assign n39594 = ~n3104 & n39593;
  assign n39595 = ~n3971 & n39594;
  assign n39596 = ~n16682 & n39595;
  assign n39597 = ~n4872 & n39596;
  assign n39598 = ~n5801 & n39597;
  assign n39599 = ~n6739 & n39598;
  assign n39600 = ~n7807 & n39599;
  assign n39601 = ~n8989 & n39600;
  assign n39602 = ~n10273 & n39601;
  assign n39603 = ~n16680 & n39602;
  assign n39604 = ~n16679 & n39603;
  assign n39605 = ~n11499 & n39604;
  assign n39606 = ~n13076 & n39605;
  assign n39607 = ~n14698 & n39606;
  assign n39608 = ~n16678 & n39607;
  assign n39609 = ~n16677 & n39608;
  assign n39610 = n16704 & n39609;
  assign n39611 = n16707 & n39610;
  assign n39612 = n16711 & n39611;
  assign n39613 = n16676 & n39612;
  assign n39614 = n16736 & n39613;
  assign n39615 = pi222 & ~n12743;
  assign n39616 = ~n12773 & n39615;
  assign n39617 = ~n12902 & n39616;
  assign n39618 = ~n17419 & n39617;
  assign n39619 = ~n17418 & n39618;
  assign n39620 = ~n14009 & n39619;
  assign n39621 = ~n16216 & n39620;
  assign n39622 = ~n16215 & n39621;
  assign n39623 = n16222 & n39622;
  assign n39624 = n17427 & n39623;
  assign n39625 = n17431 & n39624;
  assign n39626 = n16214 & n39625;
  assign n39627 = n17456 & n39626;
  assign n39628 = ~n39614 & ~n39627;
  assign n39629 = n39590 & n39628;
  assign n39630 = ~n13906 & n36403;
  assign n39631 = ~n16216 & n39630;
  assign n39632 = ~n15586 & n39631;
  assign n39633 = ~n16208 & n39632;
  assign n39634 = n17257 & n39633;
  assign n39635 = n17328 & n39634;
  assign n39636 = n17342 & n39635;
  assign n39637 = ~n13820 & n36516;
  assign n39638 = ~n16216 & n39637;
  assign n39639 = ~n14741 & n39638;
  assign n39640 = ~n16209 & n39639;
  assign n39641 = ~n16211 & n39640;
  assign n39642 = n17238 & n39641;
  assign n39643 = n17232 & n39642;
  assign n39644 = n17225 & n39643;
  assign n39645 = ~n39636 & ~n39644;
  assign n39646 = ~n14073 & n36508;
  assign n39647 = ~n16216 & n39646;
  assign n39648 = ~n15616 & n39647;
  assign n39649 = ~n16224 & n39648;
  assign n39650 = n17086 & n39649;
  assign n39651 = n17351 & n39650;
  assign n39652 = n17350 & n39651;
  assign n39653 = n17370 & n39652;
  assign n39654 = ~n13093 & n33575;
  assign n39655 = ~n16216 & n39654;
  assign n39656 = ~n16215 & n39655;
  assign n39657 = n16222 & n39656;
  assign n39658 = n17516 & n39657;
  assign n39659 = n16214 & n39658;
  assign n39660 = n17512 & n39659;
  assign n39661 = n17534 & n39660;
  assign n39662 = ~n39653 & ~n39661;
  assign n39663 = n39645 & n39662;
  assign n39664 = ~n15075 & n36425;
  assign n39665 = ~n16216 & n39664;
  assign n39666 = ~n16537 & n39665;
  assign n39667 = n16544 & n39666;
  assign n39668 = ~n16831 & n36429;
  assign n39669 = ~n16829 & n39668;
  assign n39670 = n16836 & n39669;
  assign n39671 = pi270 & ~n501;
  assign n39672 = n12872 & n39671;
  assign n39673 = n17949 & n39672;
  assign n39674 = n17954 & n39673;
  assign n39675 = n17947 & n39674;
  assign n39676 = n17982 & n39675;
  assign n39677 = ~n1172 & n39676;
  assign n39678 = ~n996 & n39677;
  assign n39679 = ~n2306 & n39678;
  assign n39680 = ~n500 & n39679;
  assign n39681 = n17940 & n39680;
  assign n39682 = n17991 & n39681;
  assign n39683 = n17938 & n39682;
  assign n39684 = n17929 & n39683;
  assign n39685 = n17921 & n39684;
  assign n39686 = n18029 & n39685;
  assign n39687 = ~n7236 & n39686;
  assign n39688 = ~n6137 & n39687;
  assign n39689 = n6193 & n39688;
  assign n39690 = n6134 & n39689;
  assign n39691 = ~n8867 & n39690;
  assign n39692 = ~n7235 & n39691;
  assign n39693 = n7296 & n39692;
  assign n39694 = n7231 & n39693;
  assign n39695 = ~n10027 & n39694;
  assign n39696 = ~n8866 & n39695;
  assign n39697 = n8898 & n39696;
  assign n39698 = n8863 & n39697;
  assign n39699 = pi278 & ~n501;
  assign n39700 = n12872 & n39699;
  assign n39701 = n18049 & n39700;
  assign n39702 = n18053 & n39701;
  assign n39703 = n18047 & n39702;
  assign n39704 = n18080 & n39703;
  assign n39705 = ~n1172 & n39704;
  assign n39706 = ~n996 & n39705;
  assign n39707 = ~n2306 & n39706;
  assign n39708 = ~n500 & n39707;
  assign n39709 = n18038 & n39708;
  assign n39710 = n18037 & n39709;
  assign n39711 = n18088 & n39710;
  assign n39712 = n18106 & n39711;
  assign n39713 = n18035 & n39712;
  assign n39714 = n18134 & n39713;
  assign n39715 = ~n7236 & n39714;
  assign n39716 = ~n6137 & n39715;
  assign n39717 = n6193 & n39716;
  assign n39718 = n6134 & n39717;
  assign n39719 = ~n8867 & n39718;
  assign n39720 = ~n7235 & n39719;
  assign n39721 = n7296 & n39720;
  assign n39722 = n7231 & n39721;
  assign n39723 = ~n10027 & n39722;
  assign n39724 = ~n8866 & n39723;
  assign n39725 = n8898 & n39724;
  assign n39726 = n8863 & n39725;
  assign n39727 = ~n39698 & ~n39726;
  assign n39728 = ~n10788 & ~n39727;
  assign n39729 = ~n10026 & n39728;
  assign n39730 = n10072 & n39729;
  assign n39731 = n10021 & n39730;
  assign n39732 = ~n39670 & ~n39731;
  assign n39733 = ~n39667 & n39732;
  assign n39734 = ~n15278 & n36500;
  assign n39735 = ~n16216 & n39734;
  assign n39736 = n16939 & n39735;
  assign n39737 = ~n16937 & n39736;
  assign n39738 = n16944 & n39737;
  assign n39739 = n16936 & n39738;
  assign n39740 = ~n15167 & n36495;
  assign n39741 = ~n16216 & n39740;
  assign n39742 = ~n16220 & n39741;
  assign n39743 = ~n16466 & n39742;
  assign n39744 = n16476 & n39743;
  assign n39745 = ~n39739 & ~n39744;
  assign n39746 = n39733 & n39745;
  assign n39747 = ~n13764 & n36410;
  assign n39748 = ~n16216 & n39747;
  assign n39749 = ~n15465 & n39748;
  assign n39750 = ~n16209 & n39749;
  assign n39751 = n17086 & n39750;
  assign n39752 = n17133 & n39751;
  assign n39753 = n17122 & n39752;
  assign n39754 = ~n13726 & n36417;
  assign n39755 = ~n16216 & n39754;
  assign n39756 = ~n15419 & n39755;
  assign n39757 = n17086 & n39756;
  assign n39758 = n17094 & n39757;
  assign n39759 = n17083 & n39758;
  assign n39760 = ~n39753 & ~n39759;
  assign n39761 = n39746 & n39760;
  assign n39762 = n39663 & n39761;
  assign n39763 = n39629 & n39762;
  assign n39764 = pi262 & ~n16417;
  assign n39765 = ~n17766 & n39764;
  assign n39766 = ~n16216 & n39765;
  assign n39767 = ~n16215 & n39766;
  assign n39768 = n16222 & n39767;
  assign n39769 = n17637 & n39768;
  assign n39770 = n17629 & n39769;
  assign n39771 = n17765 & n39770;
  assign n39772 = n17874 & n39771;
  assign n39773 = pi174 & ~n8633;
  assign n39774 = ~n8455 & n39773;
  assign n39775 = ~n8834 & n39774;
  assign n39776 = ~n10002 & n39775;
  assign n39777 = ~n17152 & n39776;
  assign n39778 = ~n17151 & n39777;
  assign n39779 = ~n11297 & n39778;
  assign n39780 = ~n12240 & n39779;
  assign n39781 = ~n13135 & n39780;
  assign n39782 = ~n16216 & n39781;
  assign n39783 = ~n16215 & n39782;
  assign n39784 = n16222 & n39783;
  assign n39785 = n17163 & n39784;
  assign n39786 = n17167 & n39785;
  assign n39787 = n17150 & n39786;
  assign n39788 = n17192 & n39787;
  assign n39789 = ~n39772 & ~n39788;
  assign n39790 = ~n6401 & n28587;
  assign n39791 = ~n6784 & n39790;
  assign n39792 = ~n7158 & n39791;
  assign n39793 = ~n8250 & n39792;
  assign n39794 = ~n9414 & n39793;
  assign n39795 = ~n16957 & n39794;
  assign n39796 = ~n16956 & n39795;
  assign n39797 = ~n10667 & n39796;
  assign n39798 = ~n12083 & n39797;
  assign n39799 = ~n13644 & n39798;
  assign n39800 = ~n16216 & n39799;
  assign n39801 = ~n16215 & n39800;
  assign n39802 = n16222 & n39801;
  assign n39803 = n16971 & n39802;
  assign n39804 = n16975 & n39803;
  assign n39805 = n16955 & n39804;
  assign n39806 = n17000 & n39805;
  assign n39807 = ~n11042 & n36376;
  assign n39808 = ~n11188 & n39807;
  assign n39809 = ~n17378 & n39808;
  assign n39810 = ~n17377 & n39809;
  assign n39811 = ~n12380 & n39810;
  assign n39812 = ~n14045 & n39811;
  assign n39813 = ~n16216 & n39812;
  assign n39814 = ~n16215 & n39813;
  assign n39815 = n16222 & n39814;
  assign n39816 = n17387 & n39815;
  assign n39817 = n17391 & n39816;
  assign n39818 = n17376 & n39817;
  assign n39819 = n17416 & n39818;
  assign n39820 = ~n39806 & ~n39819;
  assign n39821 = n39789 & n39820;
  assign n39822 = ~n9763 & n36566;
  assign n39823 = ~n9929 & n39822;
  assign n39824 = ~n17263 & n39823;
  assign n39825 = ~n17262 & n39824;
  assign n39826 = ~n11266 & n39825;
  assign n39827 = ~n11588 & n39826;
  assign n39828 = ~n13859 & n39827;
  assign n39829 = ~n16216 & n39828;
  assign n39830 = ~n16215 & n39829;
  assign n39831 = n16222 & n39830;
  assign n39832 = n17273 & n39831;
  assign n39833 = n17277 & n39832;
  assign n39834 = n17261 & n39833;
  assign n39835 = n17302 & n39834;
  assign n39836 = pi126 & ~n5686;
  assign n39837 = ~n5349 & n39836;
  assign n39838 = ~n5808 & n39837;
  assign n39839 = ~n6056 & n39838;
  assign n39840 = ~n7073 & n39839;
  assign n39841 = ~n8179 & n39840;
  assign n39842 = ~n9344 & n39841;
  assign n39843 = ~n16418 & n39842;
  assign n39844 = ~n16361 & n39843;
  assign n39845 = ~n10594 & n39844;
  assign n39846 = ~n12005 & n39845;
  assign n39847 = ~n13558 & n39846;
  assign n39848 = ~n16216 & n39847;
  assign n39849 = ~n16215 & n39848;
  assign n39850 = n16432 & n39849;
  assign n39851 = n16435 & n39850;
  assign n39852 = n16439 & n39851;
  assign n39853 = n16305 & n39852;
  assign n39854 = n16464 & n39853;
  assign n39855 = ~n39835 & ~n39854;
  assign n39856 = ~n4460 & n36582;
  assign n39857 = ~n4817 & n39856;
  assign n39858 = ~n4902 & n39857;
  assign n39859 = ~n6001 & n39858;
  assign n39860 = ~n7014 & n39859;
  assign n39861 = ~n8114 & n39860;
  assign n39862 = ~n9276 & n39861;
  assign n39863 = ~n16486 & n39862;
  assign n39864 = ~n16485 & n39863;
  assign n39865 = ~n10523 & n39864;
  assign n39866 = ~n11928 & n39865;
  assign n39867 = ~n13479 & n39866;
  assign n39868 = ~n16216 & n39867;
  assign n39869 = ~n16220 & n39868;
  assign n39870 = n16503 & n39869;
  assign n39871 = n16506 & n39870;
  assign n39872 = n16510 & n39871;
  assign n39873 = n16484 & n39872;
  assign n39874 = n16535 & n39873;
  assign n39875 = pi062 & ~n1526;
  assign n39876 = ~n1556 & n39875;
  assign n39877 = ~n2242 & n39876;
  assign n39878 = ~n3095 & n39877;
  assign n39879 = ~n3997 & n39878;
  assign n39880 = ~n4003 & n39879;
  assign n39881 = ~n4837 & n39880;
  assign n39882 = ~n5822 & n39881;
  assign n39883 = ~n6820 & n39882;
  assign n39884 = ~n7785 & n39883;
  assign n39885 = ~n9027 & n39884;
  assign n39886 = ~n10245 & n39885;
  assign n39887 = ~n16748 & n39886;
  assign n39888 = ~n16747 & n39887;
  assign n39889 = ~n11536 & n39888;
  assign n39890 = ~n13036 & n39889;
  assign n39891 = ~n14653 & n39890;
  assign n39892 = ~n16746 & n39891;
  assign n39893 = ~n16745 & n39892;
  assign n39894 = n16770 & n39893;
  assign n39895 = n16773 & n39894;
  assign n39896 = n16777 & n39895;
  assign n39897 = n16744 & n39896;
  assign n39898 = n16802 & n39897;
  assign n39899 = ~n39874 & ~n39898;
  assign n39900 = n39855 & n39899;
  assign n39901 = ~n7505 & n24592;
  assign n39902 = ~n7869 & n39901;
  assign n39903 = ~n8346 & n39902;
  assign n39904 = ~n9485 & n39903;
  assign n39905 = ~n17018 & n39904;
  assign n39906 = ~n17017 & n39905;
  assign n39907 = ~n10741 & n39906;
  assign n39908 = ~n12158 & n39907;
  assign n39909 = ~n13693 & n39908;
  assign n39910 = ~n16216 & n39909;
  assign n39911 = ~n16215 & n39910;
  assign n39912 = n16222 & n39911;
  assign n39913 = n17031 & n39912;
  assign n39914 = n17035 & n39913;
  assign n39915 = n17016 & n39914;
  assign n39916 = n17060 & n39915;
  assign n39917 = ~n16216 & n36366;
  assign n39918 = ~n16215 & n39917;
  assign n39919 = n16222 & n39918;
  assign n39920 = n16225 & n39919;
  assign n39921 = n16229 & n39920;
  assign n39922 = n16214 & n39921;
  assign n39923 = n16297 & n39922;
  assign n39924 = ~n39916 & ~n39923;
  assign n39925 = pi078 & ~n2602;
  assign n39926 = ~n2783 & n39925;
  assign n39927 = ~n3066 & n39926;
  assign n39928 = ~n3983 & n39927;
  assign n39929 = ~n4003 & n39928;
  assign n39930 = ~n4024 & n39929;
  assign n39931 = ~n4999 & n39930;
  assign n39932 = ~n5827 & n39931;
  assign n39933 = ~n6893 & n39932;
  assign n39934 = ~n7890 & n39933;
  assign n39935 = ~n9131 & n39934;
  assign n39936 = ~n16617 & n39935;
  assign n39937 = ~n16616 & n39936;
  assign n39938 = ~n10278 & n39937;
  assign n39939 = ~n11662 & n39938;
  assign n39940 = ~n13191 & n39939;
  assign n39941 = ~n16615 & n39940;
  assign n39942 = ~n16614 & n39941;
  assign n39943 = n16636 & n39942;
  assign n39944 = n16639 & n39943;
  assign n39945 = n16643 & n39944;
  assign n39946 = n16613 & n39945;
  assign n39947 = n16668 & n39946;
  assign n39948 = pi238 & ~n14350;
  assign n39949 = ~n14381 & n39948;
  assign n39950 = ~n14519 & n39949;
  assign n39951 = ~n17537 & n39950;
  assign n39952 = ~n17536 & n39951;
  assign n39953 = ~n16216 & n39952;
  assign n39954 = ~n16215 & n39953;
  assign n39955 = n16222 & n39954;
  assign n39956 = n17544 & n39955;
  assign n39957 = n17547 & n39956;
  assign n39958 = n16214 & n39957;
  assign n39959 = n17572 & n39958;
  assign n39960 = ~n39947 & ~n39959;
  assign n39961 = n39924 & n39960;
  assign n39962 = n39900 & n39961;
  assign n39963 = n39821 & n39962;
  assign po143 = ~n39763 | ~n39963;
  assign po146 = n1372 | n2242;
  assign n39966 = ~n3066 & ~n3864;
  assign po147 = n3828 | ~n39966;
  assign n39968 = ~n2242 & n3095;
  assign po148 = n3864 | n39968;
  assign n39970 = ~n3931 & ~n4002;
  assign n39971 = ~n3940 & ~n3983;
  assign po150 = ~n39970 | ~n39971;
  assign n39973 = ~n3931 & ~n3997;
  assign po151 = n3940 | ~n39973;
  assign n39975 = ~n4128 & ~n4858;
  assign po152 = n4817 | ~n39975;
  assign n39977 = n4072 & n4904;
  assign n39978 = ~n4001 & ~n4024;
  assign n39979 = ~n39977 & n39978;
  assign po153 = ~po152 & ~n39979;
  assign n39981 = ~n4001 & ~n4858;
  assign n39982 = ~n4837 & ~n39977;
  assign po154 = ~n39981 | ~n39982;
  assign n39984 = ~n4881 & ~n5769;
  assign n39985 = ~n4902 & ~n5058;
  assign n39986 = ~n5808 & n39985;
  assign po155 = ~n39984 | ~n39986;
  assign n39988 = ~n4910 & ~n4999;
  assign n39989 = ~n5043 & n39988;
  assign n39990 = ~n4881 & ~n4902;
  assign n39991 = ~n39989 & n39990;
  assign po156 = n5769 | n39991;
  assign n39993 = ~n4910 & ~n5043;
  assign n39994 = ~n5822 & n39993;
  assign n39995 = ~n4902 & ~n39994;
  assign n39996 = ~n4881 & ~n5808;
  assign po157 = n39995 | ~n39996;
  assign n39998 = ~n5967 & ~n6784;
  assign n39999 = ~n6027 & ~n6754;
  assign n40000 = n39998 & n39999;
  assign n40001 = ~n6001 & ~n6056;
  assign n40002 = ~n6114 & n40001;
  assign po158 = ~n40000 | ~n40002;
  assign n40004 = ~n5827 & n5944;
  assign n40005 = ~n6001 & ~n6027;
  assign n40006 = ~n6056 & n40005;
  assign n40007 = ~n40004 & n40006;
  assign n40008 = ~n6754 & ~n6784;
  assign n40009 = ~n6114 & n40008;
  assign po159 = n40007 | ~n40009;
  assign n40011 = n5944 & ~n6820;
  assign n40012 = ~n6001 & ~n40011;
  assign n40013 = ~n6027 & ~n6056;
  assign n40014 = ~n40012 & n40013;
  assign n40015 = ~n6114 & ~n40014;
  assign po160 = n6754 | n40015;
  assign n40017 = ~n6967 & ~n7869;
  assign n40018 = ~n7029 & ~n7095;
  assign n40019 = n40017 & n40018;
  assign n40020 = ~n7014 & ~n7073;
  assign n40021 = ~n7158 & ~n7204;
  assign n40022 = n40020 & n40021;
  assign po162 = ~n40019 | ~n40022;
  assign n40024 = ~n6893 & ~n6917;
  assign n40025 = ~n6951 & n40024;
  assign n40026 = ~n7014 & ~n7029;
  assign n40027 = ~n7073 & n40026;
  assign n40028 = ~n40025 & n40027;
  assign n40029 = ~n7095 & ~n7869;
  assign n40030 = ~n7158 & n40029;
  assign n40031 = ~n7204 & n40030;
  assign po163 = n40028 | ~n40031;
  assign n40033 = ~n6917 & ~n6951;
  assign n40034 = ~n7785 & n40033;
  assign n40035 = ~n7014 & ~n40034;
  assign n40036 = ~n7029 & ~n7073;
  assign n40037 = ~n40035 & n40036;
  assign n40038 = ~n7095 & ~n7158;
  assign n40039 = ~n40037 & n40038;
  assign n40040 = ~n7204 & ~n7869;
  assign po164 = n40039 | ~n40040;
  assign n40042 = ~n8250 & ~n8291;
  assign n40043 = ~n8346 & n40042;
  assign n40044 = ~n8053 & ~n8145;
  assign n40045 = ~n8218 & n40044;
  assign n40046 = ~n8114 & ~n8179;
  assign n40047 = n40045 & n40046;
  assign n40048 = n40043 & n40047;
  assign po166 = ~po165 & ~n40048;
  assign n40050 = ~n7890 & ~n7999;
  assign n40051 = ~n8037 & n40050;
  assign n40052 = ~n8114 & ~n8145;
  assign n40053 = ~n8179 & n40052;
  assign n40054 = ~n40051 & n40053;
  assign n40055 = ~n8218 & ~n8250;
  assign n40056 = n8347 & n40055;
  assign n40057 = ~n40054 & n40056;
  assign po167 = ~po165 & ~n40057;
  assign n40059 = ~n7999 & ~n8037;
  assign n40060 = ~n9027 & n40059;
  assign n40061 = ~n8114 & ~n40060;
  assign n40062 = ~n8145 & ~n8179;
  assign n40063 = ~n40061 & n40062;
  assign n40064 = n40055 & ~n40063;
  assign n40065 = n8347 & ~n40064;
  assign n40066 = ~n8397 & ~n40065;
  assign po168 = n8900 | n40066;
  assign n40068 = ~n9414 & ~n9453;
  assign n40069 = ~n9485 & n40068;
  assign n40070 = ~n9215 & ~n9307;
  assign n40071 = ~n9381 & n40070;
  assign n40072 = ~n9276 & ~n9344;
  assign n40073 = n40071 & n40072;
  assign n40074 = n40069 & n40073;
  assign po170 = ~po169 & ~n40074;
  assign n40076 = ~n9131 & ~n9160;
  assign n40077 = ~n9200 & n40076;
  assign n40078 = ~n9276 & ~n9307;
  assign n40079 = ~n9344 & n40078;
  assign n40080 = ~n40077 & n40079;
  assign n40081 = ~n9381 & ~n9414;
  assign n40082 = n9486 & n40081;
  assign n40083 = ~n40080 & n40082;
  assign n40084 = ~n9533 & ~n10094;
  assign n40085 = ~n10002 & n40084;
  assign n40086 = ~n40083 & n40085;
  assign po171 = n10074 | n40086;
  assign n40088 = ~n9160 & ~n9200;
  assign n40089 = ~n10245 & n40088;
  assign n40090 = ~n9276 & ~n40089;
  assign n40091 = ~n9307 & ~n9344;
  assign n40092 = ~n40090 & n40091;
  assign n40093 = n40081 & ~n40092;
  assign n40094 = n9486 & ~n40093;
  assign n40095 = ~n10002 & ~n10094;
  assign n40096 = ~n40094 & n40095;
  assign po172 = ~n9930 | n40096;
  assign n40098 = ~n10667 & ~n10705;
  assign n40099 = ~n10741 & n40098;
  assign n40100 = ~n10460 & ~n10554;
  assign n40101 = ~n10629 & n40100;
  assign n40102 = ~n10523 & ~n10594;
  assign n40103 = n40101 & n40102;
  assign n40104 = n40099 & n40103;
  assign po174 = ~po173 & ~n40104;
  assign n40106 = ~n10278 & ~n10400;
  assign n40107 = ~n10445 & n40106;
  assign n40108 = ~n10523 & ~n10554;
  assign n40109 = ~n10594 & n40108;
  assign n40110 = ~n40107 & n40109;
  assign n40111 = ~n10629 & ~n10667;
  assign n40112 = n10742 & n40111;
  assign n40113 = ~n40110 & n40112;
  assign n40114 = ~n10787 & ~n11266;
  assign n40115 = ~n11297 & ~n11318;
  assign n40116 = n40114 & n40115;
  assign n40117 = ~n40113 & n40116;
  assign n40118 = n11189 & ~n11343;
  assign po175 = n40117 | ~n40118;
  assign n40120 = ~n10400 & ~n10445;
  assign n40121 = ~n11536 & n40120;
  assign n40122 = ~n10523 & ~n40121;
  assign n40123 = ~n10554 & ~n10594;
  assign n40124 = ~n40122 & n40123;
  assign n40125 = n40111 & ~n40124;
  assign n40126 = n10742 & ~n40125;
  assign n40127 = n40115 & ~n40126;
  assign n40128 = n40114 & ~n40127;
  assign n40129 = ~n11343 & ~n40128;
  assign po176 = n10879 | n40129;
  assign n40131 = ~n12181 & ~n12240;
  assign n40132 = ~n12380 & ~n12471;
  assign n40133 = n40131 & n40132;
  assign n40134 = ~n12902 & ~n12946;
  assign n40135 = ~n11551 & n40134;
  assign n40136 = ~n11588 & ~n11611;
  assign n40137 = n40135 & n40136;
  assign po177 = ~n40133 | ~n40137;
  assign n40139 = ~n12083 & ~n12121;
  assign n40140 = ~n12158 & n40139;
  assign n40141 = ~n11860 & ~n11959;
  assign n40142 = ~n12041 & n40141;
  assign n40143 = ~n11928 & ~n12005;
  assign n40144 = n40142 & n40143;
  assign n40145 = n40140 & n40144;
  assign n40146 = ~n11551 & ~n12902;
  assign n40147 = n40136 & n40146;
  assign n40148 = n40133 & n40147;
  assign n40149 = ~n40145 & n40148;
  assign po178 = n12946 | n40149;
  assign n40151 = ~n11662 & ~n11796;
  assign n40152 = ~n11846 & n40151;
  assign n40153 = ~n11928 & ~n11959;
  assign n40154 = ~n12005 & n40153;
  assign n40155 = ~n40152 & n40154;
  assign n40156 = ~n12041 & ~n12083;
  assign n40157 = n12159 & n40156;
  assign n40158 = ~n40155 & n40157;
  assign n40159 = n40131 & n40136;
  assign n40160 = ~n40158 & n40159;
  assign n40161 = n40132 & n40146;
  assign po179 = n40160 | ~n40161;
  assign n40163 = ~n11796 & ~n11846;
  assign n40164 = ~n13036 & n40163;
  assign n40165 = ~n11928 & ~n40164;
  assign n40166 = ~n11959 & ~n12005;
  assign n40167 = ~n40165 & n40166;
  assign n40168 = n40156 & ~n40167;
  assign n40169 = n12159 & ~n40168;
  assign n40170 = n40131 & ~n40169;
  assign n40171 = n40136 & ~n40170;
  assign n40172 = ~n11551 & ~n12380;
  assign n40173 = ~n40171 & n40172;
  assign n40174 = ~n12471 & ~n12902;
  assign po180 = n40173 | ~n40174;
  assign n40176 = ~n13859 & ~n14045;
  assign n40177 = ~n14009 & ~n14073;
  assign n40178 = n40176 & n40177;
  assign n40179 = ~n14519 & ~n14568;
  assign n40180 = ~n13764 & n40179;
  assign n40181 = ~n13820 & ~n13906;
  assign n40182 = n40180 & n40181;
  assign n40183 = ~n13093 & ~n13135;
  assign n40184 = n40182 & n40183;
  assign po181 = ~n40178 | ~n40184;
  assign n40186 = ~n13407 & ~n13493;
  assign n40187 = ~n13579 & n40186;
  assign n40188 = ~n13726 & n40187;
  assign n40189 = ~n13479 & ~n13558;
  assign n40190 = ~n13644 & ~n13693;
  assign n40191 = n40189 & n40190;
  assign n40192 = n40188 & n40191;
  assign n40193 = ~n13764 & ~n13820;
  assign n40194 = ~n13906 & n40193;
  assign n40195 = ~n13135 & ~n13859;
  assign n40196 = n40194 & n40195;
  assign n40197 = n14075 & n40196;
  assign n40198 = ~n40192 & n40197;
  assign n40199 = ~n13093 & n40179;
  assign po182 = n40198 | ~n40199;
  assign n40201 = ~n13191 & ~n13318;
  assign n40202 = ~n13393 & n40201;
  assign n40203 = ~n13479 & ~n13493;
  assign n40204 = ~n13558 & n40203;
  assign n40205 = ~n40202 & n40204;
  assign n40206 = ~n13579 & ~n13726;
  assign n40207 = ~n13644 & n40206;
  assign n40208 = ~n13693 & n40207;
  assign n40209 = ~n40205 & n40208;
  assign n40210 = ~n13135 & n40193;
  assign n40211 = ~n13859 & n40210;
  assign n40212 = ~n40209 & n40211;
  assign n40213 = ~n13906 & ~n14045;
  assign n40214 = n40177 & n40213;
  assign n40215 = ~n40212 & n40214;
  assign po183 = n40199 & ~n40215;
  assign n40217 = ~n13318 & ~n13393;
  assign n40218 = ~n14653 & n40217;
  assign n40219 = ~n13479 & ~n40218;
  assign n40220 = ~n13493 & ~n13558;
  assign n40221 = ~n40219 & n40220;
  assign n40222 = ~n13579 & ~n13644;
  assign n40223 = ~n40221 & n40222;
  assign n40224 = ~n13693 & ~n13726;
  assign n40225 = ~n40223 & n40224;
  assign n40226 = ~n13135 & ~n13764;
  assign n40227 = ~n40225 & n40226;
  assign n40228 = ~n13820 & ~n13859;
  assign n40229 = ~n40227 & n40228;
  assign n40230 = n40213 & ~n40229;
  assign n40231 = n40177 & ~n40230;
  assign n40232 = ~n13093 & ~n40231;
  assign po184 = n14568 | n40232;
  assign n40234 = ~n15482 & ~n15536;
  assign n40235 = n15694 & n40234;
  assign n40236 = ~n15465 & ~n15586;
  assign n40237 = ~n15616 & n40236;
  assign n40238 = ~n16360 & ~n16417;
  assign n40239 = ~n14741 & n40238;
  assign n40240 = ~n14716 & n40239;
  assign n40241 = n15887 & n40240;
  assign n40242 = n40237 & n40241;
  assign po185 = ~n40235 | ~n40242;
  assign n40244 = ~n15075 & ~n15167;
  assign n40245 = ~n15278 & n40244;
  assign n40246 = ~n15419 & n40245;
  assign n40247 = ~n15153 & ~n15239;
  assign n40248 = ~n15330 & ~n15385;
  assign n40249 = n40247 & n40248;
  assign n40250 = n40246 & n40249;
  assign n40251 = ~n14741 & ~n15465;
  assign n40252 = n15617 & n40251;
  assign n40253 = n40235 & n40252;
  assign n40254 = ~n40250 & n40253;
  assign n40255 = ~n14716 & n40238;
  assign n40256 = n15887 & n40255;
  assign po186 = n40254 | ~n40256;
  assign n40258 = ~n14848 & ~n14980;
  assign n40259 = ~n15061 & n40258;
  assign n40260 = ~n15153 & ~n15167;
  assign n40261 = ~n15239 & n40260;
  assign n40262 = ~n40259 & n40261;
  assign n40263 = ~n15278 & ~n15419;
  assign n40264 = ~n15330 & n40263;
  assign n40265 = ~n15385 & n40264;
  assign n40266 = ~n40262 & n40265;
  assign n40267 = ~n15482 & n40251;
  assign n40268 = ~n15536 & n40267;
  assign n40269 = ~n40266 & n40268;
  assign n40270 = n15617 & ~n15657;
  assign n40271 = ~n15693 & n40270;
  assign n40272 = ~n40269 & n40271;
  assign n40273 = ~n14716 & ~n15855;
  assign n40274 = ~n15886 & n40273;
  assign n40275 = ~n40272 & n40274;
  assign po187 = n16417 | n40275;
  assign n40277 = ~n14980 & ~n15061;
  assign n40278 = ~n16255 & n40277;
  assign n40279 = ~n15153 & ~n40278;
  assign n40280 = ~n15167 & ~n15239;
  assign n40281 = ~n40279 & n40280;
  assign n40282 = ~n15278 & ~n15330;
  assign n40283 = ~n40281 & n40282;
  assign n40284 = ~n15385 & ~n15419;
  assign n40285 = ~n40283 & n40284;
  assign n40286 = ~n15465 & ~n15482;
  assign n40287 = ~n40285 & n40286;
  assign n40288 = ~n14741 & ~n15536;
  assign n40289 = ~n40287 & n40288;
  assign n40290 = ~n15586 & ~n15657;
  assign n40291 = ~n40289 & n40290;
  assign n40292 = ~n15616 & ~n15693;
  assign n40293 = ~n40291 & n40292;
  assign n40294 = n15887 & ~n40293;
  assign n40295 = ~n14716 & ~n16360;
  assign po188 = n40294 | ~n40295;
  assign n40297 = ~n17582 & ~n17737;
  assign n40298 = ~n17875 & n40297;
  assign n40299 = ~n17303 & ~n17417;
  assign n40300 = ~n17457 & ~n17573;
  assign n40301 = n40299 & n40300;
  assign n40302 = ~n17241 & ~n17343;
  assign n40303 = ~n17371 & ~n17535;
  assign n40304 = n40302 & n40303;
  assign n40305 = n12559 & n15966;
  assign n40306 = n7813 & n40305;
  assign n40307 = n14210 & n15964;
  assign n40308 = n3941 & n17944;
  assign n40309 = n40307 & n40308;
  assign n40310 = n40306 & n40309;
  assign n40311 = n14522 & n15978;
  assign n40312 = ~n751 & ~n1527;
  assign n40313 = n12562 & n40312;
  assign n40314 = n12555 & n40313;
  assign n40315 = n40311 & n40314;
  assign n40316 = n40310 & n40315;
  assign n40317 = ~n8456 & ~n14352;
  assign n40318 = ~n15989 & ~n16146;
  assign n40319 = n40317 & n40318;
  assign n40320 = ~n7328 & ~n8705;
  assign n40321 = n17959 & n40320;
  assign n40322 = n14530 & n40321;
  assign n40323 = n40319 & n40322;
  assign n40324 = n6740 & n17970;
  assign n40325 = ~n5261 & ~n5658;
  assign n40326 = n16001 & n40325;
  assign n40327 = n40324 & n40326;
  assign n40328 = n10834 & n17968;
  assign n40329 = n15986 & n40328;
  assign n40330 = n40327 & n40329;
  assign n40331 = ~n3227 & ~n3563;
  assign n40332 = n14488 & n40331;
  assign n40333 = ~n2694 & ~n3622;
  assign n40334 = n14536 & n40333;
  assign n40335 = n40332 & n40334;
  assign n40336 = n5757 & n17977;
  assign n40337 = n15997 & n40336;
  assign n40338 = n40335 & n40337;
  assign n40339 = n40330 & n40338;
  assign n40340 = n40323 & n40339;
  assign n40341 = n40316 & n40340;
  assign n40342 = ~n1172 & n40341;
  assign n40343 = ~n996 & n40342;
  assign n40344 = ~n2306 & n40343;
  assign n40345 = ~n500 & n40344;
  assign n40346 = n17940 & n40345;
  assign n40347 = n17991 & n40346;
  assign n40348 = n17938 & n40347;
  assign n40349 = n17929 & n40348;
  assign n40350 = n17921 & n40349;
  assign n40351 = n18029 & n40350;
  assign n40352 = ~n7236 & n40351;
  assign n40353 = ~n6137 & n40352;
  assign n40354 = n6193 & n40353;
  assign n40355 = n6134 & n40354;
  assign n40356 = ~n8867 & n40355;
  assign n40357 = ~n7235 & n40356;
  assign n40358 = n7296 & n40357;
  assign n40359 = n7231 & n40358;
  assign n40360 = ~n10027 & n40359;
  assign n40361 = ~n8866 & n40360;
  assign n40362 = n8898 & n40361;
  assign n40363 = n8863 & n40362;
  assign n40364 = ~n10788 & n40363;
  assign n40365 = ~n10026 & n40364;
  assign n40366 = n10072 & n40365;
  assign n40367 = n10021 & n40366;
  assign n40368 = n4798 & n15966;
  assign n40369 = n3942 & n40368;
  assign n40370 = n14194 & n18044;
  assign n40371 = n15970 & n40370;
  assign n40372 = n40369 & n40371;
  assign n40373 = n2246 & n12554;
  assign n40374 = n18049 & n40373;
  assign n40375 = n12562 & n18041;
  assign n40376 = n11407 & n40375;
  assign n40377 = n40374 & n40376;
  assign n40378 = n40372 & n40377;
  assign n40379 = ~n15989 & ~n16115;
  assign n40380 = ~n17890 & n40379;
  assign n40381 = ~n8456 & ~n14321;
  assign n40382 = n14529 & n40381;
  assign n40383 = n12904 & n18059;
  assign n40384 = n40382 & n40383;
  assign n40385 = n40380 & n40384;
  assign n40386 = n12544 & n18063;
  assign n40387 = n6741 & n40386;
  assign n40388 = n14531 & n18070;
  assign n40389 = n40387 & n40388;
  assign n40390 = ~n4373 & ~n5321;
  assign n40391 = n16363 & n40390;
  assign n40392 = n14275 & n40391;
  assign n40393 = n15997 & n16002;
  assign n40394 = n40392 & n40393;
  assign n40395 = n40389 & n40394;
  assign n40396 = n40385 & n40395;
  assign n40397 = n40378 & n40396;
  assign n40398 = ~n1172 & n40397;
  assign n40399 = ~n996 & n40398;
  assign n40400 = ~n2306 & n40399;
  assign n40401 = ~n500 & n40400;
  assign n40402 = n18038 & n40401;
  assign n40403 = n18037 & n40402;
  assign n40404 = n18088 & n40403;
  assign n40405 = n18106 & n40404;
  assign n40406 = n18035 & n40405;
  assign n40407 = n18134 & n40406;
  assign n40408 = ~n7236 & n40407;
  assign n40409 = ~n6137 & n40408;
  assign n40410 = n6193 & n40409;
  assign n40411 = n6134 & n40410;
  assign n40412 = ~n8867 & n40411;
  assign n40413 = ~n7235 & n40412;
  assign n40414 = n7296 & n40413;
  assign n40415 = n7231 & n40414;
  assign n40416 = ~n10027 & n40415;
  assign n40417 = ~n8866 & n40416;
  assign n40418 = n8898 & n40417;
  assign n40419 = n8863 & n40418;
  assign n40420 = ~n10788 & n40419;
  assign n40421 = ~n10026 & n40420;
  assign n40422 = n10072 & n40421;
  assign n40423 = n10021 & n40422;
  assign n40424 = ~n40367 & ~n40423;
  assign n40425 = ~n17135 & n40424;
  assign n40426 = ~n17193 & n40425;
  assign n40427 = n40304 & n40426;
  assign n40428 = n40301 & n40427;
  assign po189 = ~n40298 | ~n40428;
  assign n40430 = ~n16477 & ~n16545;
  assign n40431 = ~n16946 & n40430;
  assign n40432 = ~n17096 & n40431;
  assign n40433 = ~n16465 & ~n16536;
  assign n40434 = ~n17001 & ~n17061;
  assign n40435 = n40433 & n40434;
  assign n40436 = n40432 & n40435;
  assign n40437 = ~n17135 & ~n17241;
  assign n40438 = n17372 & n40437;
  assign n40439 = ~n17193 & ~n17303;
  assign n40440 = n17458 & n40439;
  assign n40441 = n40438 & n40440;
  assign n40442 = ~n40436 & n40441;
  assign n40443 = ~n17535 & n40424;
  assign n40444 = ~n17573 & n40443;
  assign n40445 = n40298 & n40444;
  assign po190 = n40442 | ~n40445;
  assign n40447 = ~n16669 & ~n16837;
  assign n40448 = ~n16859 & n40447;
  assign n40449 = ~n16465 & ~n16477;
  assign n40450 = ~n16536 & n40449;
  assign n40451 = ~n40448 & n40450;
  assign n40452 = ~n16946 & ~n17096;
  assign n40453 = ~n17001 & n40452;
  assign n40454 = ~n17061 & n40453;
  assign n40455 = ~n40451 & n40454;
  assign n40456 = ~n17193 & n40437;
  assign n40457 = ~n17303 & n40456;
  assign n40458 = ~n40455 & n40457;
  assign n40459 = n17372 & ~n17417;
  assign n40460 = ~n17457 & n40459;
  assign n40461 = ~n40458 & n40460;
  assign n40462 = n17574 & n40297;
  assign n40463 = ~n40461 & n40462;
  assign n40464 = ~n17875 & n40424;
  assign po191 = n40463 | ~n40464;
  assign n40466 = n1557 & ~n2242;
  assign n40467 = ~n3095 & n40466;
  assign n40468 = ~n3997 & n40467;
  assign n40469 = ~n4003 & n40468;
  assign n40470 = ~n4837 & n40469;
  assign n40471 = ~n5822 & n40470;
  assign n40472 = ~n6820 & n40471;
  assign n40473 = ~n7785 & n40472;
  assign n40474 = ~n9027 & n40473;
  assign n40475 = ~n10245 & n40474;
  assign n40476 = ~n16748 & n40475;
  assign n40477 = ~n16747 & n40476;
  assign n40478 = ~n11536 & n40477;
  assign n40479 = ~n13036 & n40478;
  assign n40480 = ~n14653 & n40479;
  assign n40481 = ~n16746 & n40480;
  assign n40482 = ~n16745 & n40481;
  assign n40483 = n16770 & n40482;
  assign n40484 = n16773 & n40483;
  assign n40485 = n16777 & n40484;
  assign n40486 = n16744 & n40485;
  assign n40487 = n16802 & n40486;
  assign n40488 = ~n16837 & ~n16859;
  assign n40489 = ~n40487 & n40488;
  assign n40490 = ~n16536 & ~n40489;
  assign n40491 = n40449 & ~n40490;
  assign n40492 = ~n16946 & ~n17001;
  assign n40493 = ~n40491 & n40492;
  assign n40494 = ~n17061 & ~n17096;
  assign n40495 = ~n40493 & n40494;
  assign n40496 = ~n17135 & ~n17193;
  assign n40497 = ~n40495 & n40496;
  assign n40498 = ~n17241 & ~n17303;
  assign n40499 = ~n40497 & n40498;
  assign n40500 = ~n17343 & ~n17417;
  assign n40501 = ~n40499 & n40500;
  assign n40502 = ~n17371 & ~n17457;
  assign n40503 = ~n40501 & n40502;
  assign n40504 = n17574 & ~n40503;
  assign n40505 = n40297 & ~n40504;
  assign n40506 = ~n17875 & ~n40505;
  assign po192 = n40423 | n40506;
  assign po000 = pi000;
  assign po016 = pi031;
  assign po017 = pi032;
  assign po018 = pi033;
  assign po019 = pi034;
  assign po020 = pi035;
  assign po021 = pi036;
  assign po022 = pi037;
  assign po023 = pi038;
endmodule


